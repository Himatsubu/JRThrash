/*
TimeStamp:	2016/10/12		16:46
*/


module P3_2dim(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 8:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 5:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 5:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [14:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [14:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [14:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [14:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [14:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [14:0] w_fld_V_3_addr_0;
	wire        [31:0] w_fld_V_3_datain_0;
	wire        [31:0] w_fld_V_3_dataout_0;
	wire               w_fld_V_3_r_w_0;
	wire               w_fld_V_3_ce_0;
	reg  signed [14:0] r_fld_V_3_addr_1;
	reg         [31:0] r_fld_V_3_datain_1;
	wire        [31:0] w_fld_V_3_dataout_1;
	reg                r_fld_V_3_r_w_1;
	wire               w_fld_V_3_ce_1;
	reg  signed [31:0] r_run_k_20;
	reg  signed [31:0] r_run_j_21;
	reg  signed [31:0] r_run_n_22;
	reg  signed [31:0] r_run_mx_23;
	reg  signed [31:0] r_run_my_24;
	reg         [31:0] r_run_dt_25;
	reg         [31:0] r_run_dx_26;
	reg         [31:0] r_run_dy_27;
	reg         [31:0] r_run_r1_28;
	reg         [31:0] r_run_r2_29;
	reg         [31:0] r_run_r3_30;
	reg         [31:0] r_run_r4_31;
	reg         [31:0] r_run_YY_32;
	reg  signed [31:0] r_run_kx_33;
	reg  signed [31:0] r_run_ky_34;
	reg  signed [31:0] r_run_nlast_35;
	reg  signed [31:0] r_run_copy0_j_36;
	reg  signed [31:0] r_run_copy1_j_37;
	reg  signed [31:0] r_run_copy2_j_38;
	reg  signed [31:0] r_run_copy0_j_39;
	reg  signed [31:0] r_run_copy1_j_40;
	reg  signed [31:0] r_run_copy2_j_41;
	reg  signed [31:0] r_run_copy3_j_42;
	reg  signed [31:0] r_run_copy4_j_43;
	reg  signed [31:0] r_run_copy0_j_44;
	reg  signed [31:0] r_run_copy1_j_45;
	reg  signed [31:0] r_run_copy2_j_46;
	reg  signed [31:0] r_run_copy3_j_47;
	reg  signed [31:0] r_run_copy4_j_48;
	reg  signed [31:0] r_run_copy0_j_49;
	reg  signed [31:0] r_run_copy1_j_50;
	reg  signed [31:0] r_run_copy2_j_51;
	reg  signed [31:0] r_run_copy3_j_52;
	reg  signed [31:0] r_run_copy4_j_53;
	reg  signed [31:0] r_run_copy0_j_54;
	reg  signed [31:0] r_run_copy1_j_55;
	reg  signed [31:0] r_run_copy2_j_56;
	reg  signed [31:0] r_run_copy3_j_57;
	reg  signed [31:0] r_run_copy4_j_58;
	reg  signed [31:0] r_run_copy0_j_59;
	reg  signed [31:0] r_run_copy1_j_60;
	reg  signed [31:0] r_run_copy2_j_61;
	reg  signed [31:0] r_run_copy3_j_62;
	reg  signed [31:0] r_run_copy4_j_63;
	reg  signed [31:0] r_run_copy0_j_64;
	reg  signed [31:0] r_run_copy1_j_65;
	reg  signed [31:0] r_run_copy2_j_66;
	reg  signed [31:0] r_run_copy3_j_67;
	reg  signed [31:0] r_run_copy4_j_68;
	reg  signed [31:0] r_run_copy0_j_69;
	reg  signed [31:0] r_run_copy1_j_70;
	reg  signed [31:0] r_run_copy2_j_71;
	reg  signed [31:0] r_run_copy3_j_72;
	reg  signed [31:0] r_run_copy4_j_73;
	reg  signed [31:0] r_run_copy0_j_74;
	reg  signed [31:0] r_run_copy1_j_75;
	reg  signed [31:0] r_run_copy2_j_76;
	reg  signed [31:0] r_run_copy3_j_77;
	reg  signed [31:0] r_run_copy4_j_78;
	reg  signed [31:0] r_run_copy0_j_79;
	reg  signed [31:0] r_run_copy1_j_80;
	reg  signed [31:0] r_run_copy2_j_81;
	reg  signed [31:0] r_run_copy3_j_82;
	reg  signed [31:0] r_run_copy4_j_83;
	reg  signed [31:0] r_run_copy0_j_84;
	reg  signed [31:0] r_run_copy1_j_85;
	reg  signed [31:0] r_run_copy2_j_86;
	reg  signed [31:0] r_run_copy3_j_87;
	reg  signed [31:0] r_run_copy4_j_88;
	reg  signed [31:0] r_run_copy0_j_89;
	reg  signed [31:0] r_run_copy1_j_90;
	reg  signed [31:0] r_run_copy2_j_91;
	reg  signed [31:0] r_run_copy3_j_92;
	reg  signed [31:0] r_run_copy4_j_93;
	reg  signed [31:0] r_run_copy0_j_94;
	reg  signed [31:0] r_run_copy1_j_95;
	reg  signed [31:0] r_run_copy2_j_96;
	reg  signed [31:0] r_run_copy3_j_97;
	reg  signed [31:0] r_run_copy4_j_98;
	reg  signed [31:0] r_run_copy0_j_99;
	reg  signed [31:0] r_run_copy1_j_100;
	reg  signed [31:0] r_run_copy2_j_101;
	reg  signed [31:0] r_run_copy3_j_102;
	reg  signed [31:0] r_run_copy4_j_103;
	reg  signed [31:0] r_run_copy0_j_104;
	reg  signed [31:0] r_run_copy1_j_105;
	reg  signed [31:0] r_run_copy2_j_106;
	reg  signed [31:0] r_run_copy3_j_107;
	reg  signed [31:0] r_run_copy4_j_108;
	reg  signed [31:0] r_run_copy0_j_109;
	reg  signed [31:0] r_run_copy1_j_110;
	reg  signed [31:0] r_run_copy2_j_111;
	reg  signed [31:0] r_run_copy3_j_112;
	reg  signed [31:0] r_run_copy4_j_113;
	reg  signed [31:0] r_run_copy0_j_114;
	reg  signed [31:0] r_run_copy1_j_115;
	reg  signed [31:0] r_run_copy2_j_116;
	reg  signed [31:0] r_run_copy3_j_117;
	reg  signed [31:0] r_run_copy4_j_118;
	reg  signed [31:0] r_run_copy0_j_119;
	reg  signed [31:0] r_run_copy1_j_120;
	reg  signed [31:0] r_run_copy2_j_121;
	reg  signed [31:0] r_run_copy3_j_122;
	reg  signed [31:0] r_run_copy4_j_123;
	reg  signed [31:0] r_run_copy5_j_124;
	reg  signed [31:0] r_run_copy6_j_125;
	reg  signed [31:0] r_run_copy7_j_126;
	reg  signed [31:0] r_run_copy8_j_127;
	reg  signed [31:0] r_run_copy9_j_128;
	reg  signed [31:0] r_run_copy10_j_129;
	reg  signed [31:0] r_run_copy0_j_130;
	reg  signed [31:0] r_run_copy1_j_131;
	reg  signed [31:0] r_run_copy2_j_132;
	reg  signed [31:0] r_run_copy3_j_133;
	reg  signed [31:0] r_run_copy4_j_134;
	reg  signed [31:0] r_run_copy5_j_135;
	reg  signed [31:0] r_run_copy6_j_136;
	reg  signed [31:0] r_run_copy7_j_137;
	reg  signed [31:0] r_run_copy8_j_138;
	reg  signed [31:0] r_run_copy9_j_139;
	reg  signed [31:0] r_run_copy10_j_140;
	reg  signed [31:0] r_run_copy0_j_141;
	reg  signed [31:0] r_run_copy1_j_142;
	reg  signed [31:0] r_run_copy2_j_143;
	reg  signed [31:0] r_run_copy3_j_144;
	reg  signed [31:0] r_run_copy4_j_145;
	reg  signed [31:0] r_run_copy5_j_146;
	reg  signed [31:0] r_run_copy6_j_147;
	reg  signed [31:0] r_run_copy7_j_148;
	reg  signed [31:0] r_run_copy8_j_149;
	reg  signed [31:0] r_run_copy9_j_150;
	reg  signed [31:0] r_run_copy10_j_151;
	reg  signed [31:0] r_run_copy0_j_152;
	reg  signed [31:0] r_run_copy1_j_153;
	reg  signed [31:0] r_run_copy2_j_154;
	reg  signed [31:0] r_run_copy3_j_155;
	reg  signed [31:0] r_run_copy4_j_156;
	reg  signed [31:0] r_run_copy5_j_157;
	reg  signed [31:0] r_run_copy6_j_158;
	reg  signed [31:0] r_run_copy7_j_159;
	reg  signed [31:0] r_run_copy8_j_160;
	reg  signed [31:0] r_run_copy9_j_161;
	reg  signed [31:0] r_run_copy10_j_162;
	reg  signed [31:0] r_run_copy0_j_163;
	reg  signed [31:0] r_run_copy0_j_164;
	reg  signed [31:0] r_run_copy0_j_165;
	reg  signed [31:0] r_run_copy0_j_166;
	reg  signed [31:0] r_run_copy0_j_167;
	reg  signed [31:0] r_run_copy0_j_168;
	reg  signed [31:0] r_run_copy0_j_169;
	reg  signed [31:0] r_run_copy0_j_170;
	reg  signed [31:0] r_run_copy0_j_171;
	reg  signed [31:0] r_run_copy0_j_172;
	reg  signed [31:0] r_run_copy0_j_173;
	reg  signed [31:0] r_run_copy0_j_174;
	reg  signed [31:0] r_run_copy0_j_175;
	reg  signed [31:0] r_run_copy0_j_176;
	reg  signed [31:0] r_run_copy0_j_177;
	reg  signed [31:0] r_run_copy0_j_178;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [14:0] w_sub09_T_addr;
	reg  signed [14:0] r_sub09_T_addr;
	wire        [31:0] w_sub09_T_datain;
	reg         [31:0] r_sub09_T_datain;
	wire        [31:0] w_sub09_T_dataout;
	wire               w_sub09_T_r_w;
	reg                r_sub09_T_r_w;
	wire signed [14:0] w_sub09_V_addr;
	reg  signed [14:0] r_sub09_V_addr;
	wire        [31:0] w_sub09_V_datain;
	reg         [31:0] r_sub09_V_datain;
	wire        [31:0] w_sub09_V_dataout;
	wire               w_sub09_V_r_w;
	reg                r_sub09_V_r_w;
	wire signed [14:0] w_sub09_U_addr;
	reg  signed [14:0] r_sub09_U_addr;
	wire        [31:0] w_sub09_U_datain;
	reg         [31:0] r_sub09_U_datain;
	wire        [31:0] w_sub09_U_dataout;
	wire               w_sub09_U_r_w;
	reg                r_sub09_U_r_w;
	wire signed [14:0] w_sub09_result_addr;
	reg  signed [14:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [14:0] w_sub08_T_addr;
	reg  signed [14:0] r_sub08_T_addr;
	wire        [31:0] w_sub08_T_datain;
	reg         [31:0] r_sub08_T_datain;
	wire        [31:0] w_sub08_T_dataout;
	wire               w_sub08_T_r_w;
	reg                r_sub08_T_r_w;
	wire signed [14:0] w_sub08_V_addr;
	reg  signed [14:0] r_sub08_V_addr;
	wire        [31:0] w_sub08_V_datain;
	reg         [31:0] r_sub08_V_datain;
	wire        [31:0] w_sub08_V_dataout;
	wire               w_sub08_V_r_w;
	reg                r_sub08_V_r_w;
	wire signed [14:0] w_sub08_U_addr;
	reg  signed [14:0] r_sub08_U_addr;
	wire        [31:0] w_sub08_U_datain;
	reg         [31:0] r_sub08_U_datain;
	wire        [31:0] w_sub08_U_dataout;
	wire               w_sub08_U_r_w;
	reg                r_sub08_U_r_w;
	wire signed [14:0] w_sub08_result_addr;
	reg  signed [14:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [14:0] w_sub12_T_addr;
	reg  signed [14:0] r_sub12_T_addr;
	wire        [31:0] w_sub12_T_datain;
	reg         [31:0] r_sub12_T_datain;
	wire        [31:0] w_sub12_T_dataout;
	wire               w_sub12_T_r_w;
	reg                r_sub12_T_r_w;
	wire signed [14:0] w_sub12_V_addr;
	reg  signed [14:0] r_sub12_V_addr;
	wire        [31:0] w_sub12_V_datain;
	reg         [31:0] r_sub12_V_datain;
	wire        [31:0] w_sub12_V_dataout;
	wire               w_sub12_V_r_w;
	reg                r_sub12_V_r_w;
	wire signed [14:0] w_sub12_U_addr;
	reg  signed [14:0] r_sub12_U_addr;
	wire        [31:0] w_sub12_U_datain;
	reg         [31:0] r_sub12_U_datain;
	wire        [31:0] w_sub12_U_dataout;
	wire               w_sub12_U_r_w;
	reg                r_sub12_U_r_w;
	wire signed [14:0] w_sub12_result_addr;
	reg  signed [14:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [14:0] w_sub03_T_addr;
	reg  signed [14:0] r_sub03_T_addr;
	wire        [31:0] w_sub03_T_datain;
	reg         [31:0] r_sub03_T_datain;
	wire        [31:0] w_sub03_T_dataout;
	wire               w_sub03_T_r_w;
	reg                r_sub03_T_r_w;
	wire signed [14:0] w_sub03_V_addr;
	reg  signed [14:0] r_sub03_V_addr;
	wire        [31:0] w_sub03_V_datain;
	reg         [31:0] r_sub03_V_datain;
	wire        [31:0] w_sub03_V_dataout;
	wire               w_sub03_V_r_w;
	reg                r_sub03_V_r_w;
	wire signed [14:0] w_sub03_U_addr;
	reg  signed [14:0] r_sub03_U_addr;
	wire        [31:0] w_sub03_U_datain;
	reg         [31:0] r_sub03_U_datain;
	wire        [31:0] w_sub03_U_dataout;
	wire               w_sub03_U_r_w;
	reg                r_sub03_U_r_w;
	wire signed [14:0] w_sub03_result_addr;
	reg  signed [14:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [14:0] w_sub02_T_addr;
	reg  signed [14:0] r_sub02_T_addr;
	wire        [31:0] w_sub02_T_datain;
	reg         [31:0] r_sub02_T_datain;
	wire        [31:0] w_sub02_T_dataout;
	wire               w_sub02_T_r_w;
	reg                r_sub02_T_r_w;
	wire signed [14:0] w_sub02_V_addr;
	reg  signed [14:0] r_sub02_V_addr;
	wire        [31:0] w_sub02_V_datain;
	reg         [31:0] r_sub02_V_datain;
	wire        [31:0] w_sub02_V_dataout;
	wire               w_sub02_V_r_w;
	reg                r_sub02_V_r_w;
	wire signed [14:0] w_sub02_U_addr;
	reg  signed [14:0] r_sub02_U_addr;
	wire        [31:0] w_sub02_U_datain;
	reg         [31:0] r_sub02_U_datain;
	wire        [31:0] w_sub02_U_dataout;
	wire               w_sub02_U_r_w;
	reg                r_sub02_U_r_w;
	wire signed [14:0] w_sub02_result_addr;
	reg  signed [14:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [14:0] w_sub11_T_addr;
	reg  signed [14:0] r_sub11_T_addr;
	wire        [31:0] w_sub11_T_datain;
	reg         [31:0] r_sub11_T_datain;
	wire        [31:0] w_sub11_T_dataout;
	wire               w_sub11_T_r_w;
	reg                r_sub11_T_r_w;
	wire signed [14:0] w_sub11_V_addr;
	reg  signed [14:0] r_sub11_V_addr;
	wire        [31:0] w_sub11_V_datain;
	reg         [31:0] r_sub11_V_datain;
	wire        [31:0] w_sub11_V_dataout;
	wire               w_sub11_V_r_w;
	reg                r_sub11_V_r_w;
	wire signed [14:0] w_sub11_U_addr;
	reg  signed [14:0] r_sub11_U_addr;
	wire        [31:0] w_sub11_U_datain;
	reg         [31:0] r_sub11_U_datain;
	wire        [31:0] w_sub11_U_dataout;
	wire               w_sub11_U_r_w;
	reg                r_sub11_U_r_w;
	wire signed [14:0] w_sub11_result_addr;
	reg  signed [14:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [14:0] w_sub14_T_addr;
	reg  signed [14:0] r_sub14_T_addr;
	wire        [31:0] w_sub14_T_datain;
	reg         [31:0] r_sub14_T_datain;
	wire        [31:0] w_sub14_T_dataout;
	wire               w_sub14_T_r_w;
	reg                r_sub14_T_r_w;
	wire signed [14:0] w_sub14_V_addr;
	reg  signed [14:0] r_sub14_V_addr;
	wire        [31:0] w_sub14_V_datain;
	reg         [31:0] r_sub14_V_datain;
	wire        [31:0] w_sub14_V_dataout;
	wire               w_sub14_V_r_w;
	reg                r_sub14_V_r_w;
	wire signed [14:0] w_sub14_U_addr;
	reg  signed [14:0] r_sub14_U_addr;
	wire        [31:0] w_sub14_U_datain;
	reg         [31:0] r_sub14_U_datain;
	wire        [31:0] w_sub14_U_dataout;
	wire               w_sub14_U_r_w;
	reg                r_sub14_U_r_w;
	wire signed [14:0] w_sub14_result_addr;
	reg  signed [14:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [14:0] w_sub01_T_addr;
	reg  signed [14:0] r_sub01_T_addr;
	wire        [31:0] w_sub01_T_datain;
	reg         [31:0] r_sub01_T_datain;
	wire        [31:0] w_sub01_T_dataout;
	wire               w_sub01_T_r_w;
	reg                r_sub01_T_r_w;
	wire signed [14:0] w_sub01_V_addr;
	reg  signed [14:0] r_sub01_V_addr;
	wire        [31:0] w_sub01_V_datain;
	reg         [31:0] r_sub01_V_datain;
	wire        [31:0] w_sub01_V_dataout;
	wire               w_sub01_V_r_w;
	reg                r_sub01_V_r_w;
	wire signed [14:0] w_sub01_U_addr;
	reg  signed [14:0] r_sub01_U_addr;
	wire        [31:0] w_sub01_U_datain;
	reg         [31:0] r_sub01_U_datain;
	wire        [31:0] w_sub01_U_dataout;
	wire               w_sub01_U_r_w;
	reg                r_sub01_U_r_w;
	wire signed [14:0] w_sub01_result_addr;
	reg  signed [14:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [14:0] w_sub13_T_addr;
	reg  signed [14:0] r_sub13_T_addr;
	wire        [31:0] w_sub13_T_datain;
	reg         [31:0] r_sub13_T_datain;
	wire        [31:0] w_sub13_T_dataout;
	wire               w_sub13_T_r_w;
	reg                r_sub13_T_r_w;
	wire signed [14:0] w_sub13_V_addr;
	reg  signed [14:0] r_sub13_V_addr;
	wire        [31:0] w_sub13_V_datain;
	reg         [31:0] r_sub13_V_datain;
	wire        [31:0] w_sub13_V_dataout;
	wire               w_sub13_V_r_w;
	reg                r_sub13_V_r_w;
	wire signed [14:0] w_sub13_U_addr;
	reg  signed [14:0] r_sub13_U_addr;
	wire        [31:0] w_sub13_U_datain;
	reg         [31:0] r_sub13_U_datain;
	wire        [31:0] w_sub13_U_dataout;
	wire               w_sub13_U_r_w;
	reg                r_sub13_U_r_w;
	wire signed [14:0] w_sub13_result_addr;
	reg  signed [14:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [14:0] w_sub00_T_addr;
	reg  signed [14:0] r_sub00_T_addr;
	wire        [31:0] w_sub00_T_datain;
	reg         [31:0] r_sub00_T_datain;
	wire        [31:0] w_sub00_T_dataout;
	wire               w_sub00_T_r_w;
	reg                r_sub00_T_r_w;
	wire signed [14:0] w_sub00_V_addr;
	reg  signed [14:0] r_sub00_V_addr;
	wire        [31:0] w_sub00_V_datain;
	reg         [31:0] r_sub00_V_datain;
	wire        [31:0] w_sub00_V_dataout;
	wire               w_sub00_V_r_w;
	reg                r_sub00_V_r_w;
	wire signed [14:0] w_sub00_U_addr;
	reg  signed [14:0] r_sub00_U_addr;
	wire        [31:0] w_sub00_U_datain;
	reg         [31:0] r_sub00_U_datain;
	wire        [31:0] w_sub00_U_dataout;
	wire               w_sub00_U_r_w;
	reg                r_sub00_U_r_w;
	wire signed [14:0] w_sub00_result_addr;
	reg  signed [14:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [14:0] w_sub07_T_addr;
	reg  signed [14:0] r_sub07_T_addr;
	wire        [31:0] w_sub07_T_datain;
	reg         [31:0] r_sub07_T_datain;
	wire        [31:0] w_sub07_T_dataout;
	wire               w_sub07_T_r_w;
	reg                r_sub07_T_r_w;
	wire signed [14:0] w_sub07_V_addr;
	reg  signed [14:0] r_sub07_V_addr;
	wire        [31:0] w_sub07_V_datain;
	reg         [31:0] r_sub07_V_datain;
	wire        [31:0] w_sub07_V_dataout;
	wire               w_sub07_V_r_w;
	reg                r_sub07_V_r_w;
	wire signed [14:0] w_sub07_U_addr;
	reg  signed [14:0] r_sub07_U_addr;
	wire        [31:0] w_sub07_U_datain;
	reg         [31:0] r_sub07_U_datain;
	wire        [31:0] w_sub07_U_dataout;
	wire               w_sub07_U_r_w;
	reg                r_sub07_U_r_w;
	wire signed [14:0] w_sub07_result_addr;
	reg  signed [14:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [14:0] w_sub06_T_addr;
	reg  signed [14:0] r_sub06_T_addr;
	wire        [31:0] w_sub06_T_datain;
	reg         [31:0] r_sub06_T_datain;
	wire        [31:0] w_sub06_T_dataout;
	wire               w_sub06_T_r_w;
	reg                r_sub06_T_r_w;
	wire signed [14:0] w_sub06_V_addr;
	reg  signed [14:0] r_sub06_V_addr;
	wire        [31:0] w_sub06_V_datain;
	reg         [31:0] r_sub06_V_datain;
	wire        [31:0] w_sub06_V_dataout;
	wire               w_sub06_V_r_w;
	reg                r_sub06_V_r_w;
	wire signed [14:0] w_sub06_U_addr;
	reg  signed [14:0] r_sub06_U_addr;
	wire        [31:0] w_sub06_U_datain;
	reg         [31:0] r_sub06_U_datain;
	wire        [31:0] w_sub06_U_dataout;
	wire               w_sub06_U_r_w;
	reg                r_sub06_U_r_w;
	wire signed [14:0] w_sub06_result_addr;
	reg  signed [14:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [14:0] w_sub15_T_addr;
	reg  signed [14:0] r_sub15_T_addr;
	wire        [31:0] w_sub15_T_datain;
	reg         [31:0] r_sub15_T_datain;
	wire        [31:0] w_sub15_T_dataout;
	wire               w_sub15_T_r_w;
	reg                r_sub15_T_r_w;
	wire signed [14:0] w_sub15_V_addr;
	reg  signed [14:0] r_sub15_V_addr;
	wire        [31:0] w_sub15_V_datain;
	reg         [31:0] r_sub15_V_datain;
	wire        [31:0] w_sub15_V_dataout;
	wire               w_sub15_V_r_w;
	reg                r_sub15_V_r_w;
	wire signed [14:0] w_sub15_U_addr;
	reg  signed [14:0] r_sub15_U_addr;
	wire        [31:0] w_sub15_U_datain;
	reg         [31:0] r_sub15_U_datain;
	wire        [31:0] w_sub15_U_dataout;
	wire               w_sub15_U_r_w;
	reg                r_sub15_U_r_w;
	wire signed [14:0] w_sub15_result_addr;
	reg  signed [14:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [14:0] w_sub05_T_addr;
	reg  signed [14:0] r_sub05_T_addr;
	wire        [31:0] w_sub05_T_datain;
	reg         [31:0] r_sub05_T_datain;
	wire        [31:0] w_sub05_T_dataout;
	wire               w_sub05_T_r_w;
	reg                r_sub05_T_r_w;
	wire signed [14:0] w_sub05_V_addr;
	reg  signed [14:0] r_sub05_V_addr;
	wire        [31:0] w_sub05_V_datain;
	reg         [31:0] r_sub05_V_datain;
	wire        [31:0] w_sub05_V_dataout;
	wire               w_sub05_V_r_w;
	reg                r_sub05_V_r_w;
	wire signed [14:0] w_sub05_U_addr;
	reg  signed [14:0] r_sub05_U_addr;
	wire        [31:0] w_sub05_U_datain;
	reg         [31:0] r_sub05_U_datain;
	wire        [31:0] w_sub05_U_dataout;
	wire               w_sub05_U_r_w;
	reg                r_sub05_U_r_w;
	wire signed [14:0] w_sub05_result_addr;
	reg  signed [14:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [14:0] w_sub04_T_addr;
	reg  signed [14:0] r_sub04_T_addr;
	wire        [31:0] w_sub04_T_datain;
	reg         [31:0] r_sub04_T_datain;
	wire        [31:0] w_sub04_T_dataout;
	wire               w_sub04_T_r_w;
	reg                r_sub04_T_r_w;
	wire signed [14:0] w_sub04_V_addr;
	reg  signed [14:0] r_sub04_V_addr;
	wire        [31:0] w_sub04_V_datain;
	reg         [31:0] r_sub04_V_datain;
	wire        [31:0] w_sub04_V_dataout;
	wire               w_sub04_V_r_w;
	reg                r_sub04_V_r_w;
	wire signed [14:0] w_sub04_U_addr;
	reg  signed [14:0] r_sub04_U_addr;
	wire        [31:0] w_sub04_U_datain;
	reg         [31:0] r_sub04_U_datain;
	wire        [31:0] w_sub04_U_dataout;
	wire               w_sub04_U_r_w;
	reg                r_sub04_U_r_w;
	wire signed [14:0] w_sub04_result_addr;
	reg  signed [14:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [14:0] w_sub10_T_addr;
	reg  signed [14:0] r_sub10_T_addr;
	wire        [31:0] w_sub10_T_datain;
	reg         [31:0] r_sub10_T_datain;
	wire        [31:0] w_sub10_T_dataout;
	wire               w_sub10_T_r_w;
	reg                r_sub10_T_r_w;
	wire signed [14:0] w_sub10_V_addr;
	reg  signed [14:0] r_sub10_V_addr;
	wire        [31:0] w_sub10_V_datain;
	reg         [31:0] r_sub10_V_datain;
	wire        [31:0] w_sub10_V_dataout;
	wire               w_sub10_V_r_w;
	reg                r_sub10_V_r_w;
	wire signed [14:0] w_sub10_U_addr;
	reg  signed [14:0] r_sub10_U_addr;
	wire        [31:0] w_sub10_U_datain;
	reg         [31:0] r_sub10_U_datain;
	wire        [31:0] w_sub10_U_dataout;
	wire               w_sub10_U_r_w;
	reg                r_sub10_U_r_w;
	wire signed [14:0] w_sub10_result_addr;
	reg  signed [14:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire               w_sys_tmp12;
	wire               w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp15;
	wire               w_sys_tmp16;
	wire        [31:0] w_sys_tmp18;
	wire        [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire        [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp27;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp32;
	wire signed [31:0] w_sys_tmp33;
	wire        [31:0] w_sys_tmp36;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp45;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire        [31:0] w_sys_tmp128;
	wire               w_sys_tmp226;
	wire               w_sys_tmp227;
	wire signed [31:0] w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire               w_sys_tmp230;
	wire               w_sys_tmp231;
	wire signed [31:0] w_sys_tmp232;
	wire signed [31:0] w_sys_tmp235;
	wire signed [31:0] w_sys_tmp236;
	wire signed [31:0] w_sys_tmp237;
	wire        [31:0] w_sys_tmp238;
	wire signed [31:0] w_sys_tmp239;
	wire signed [31:0] w_sys_tmp240;
	wire signed [31:0] w_sys_tmp243;
	wire signed [31:0] w_sys_tmp244;
	wire        [31:0] w_sys_tmp246;
	wire signed [31:0] w_sys_tmp247;
	wire signed [31:0] w_sys_tmp248;
	wire signed [31:0] w_sys_tmp251;
	wire signed [31:0] w_sys_tmp252;
	wire        [31:0] w_sys_tmp254;
	wire signed [31:0] w_sys_tmp255;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp258;
	wire signed [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp260;
	wire signed [31:0] w_sys_tmp261;
	wire signed [31:0] w_sys_tmp262;
	wire signed [31:0] w_sys_tmp263;
	wire signed [31:0] w_sys_tmp444;
	wire               w_sys_tmp445;
	wire               w_sys_tmp446;
	wire signed [31:0] w_sys_tmp447;
	wire signed [31:0] w_sys_tmp450;
	wire signed [31:0] w_sys_tmp451;
	wire signed [31:0] w_sys_tmp452;
	wire        [31:0] w_sys_tmp453;
	wire signed [31:0] w_sys_tmp454;
	wire signed [31:0] w_sys_tmp455;
	wire signed [31:0] w_sys_tmp458;
	wire signed [31:0] w_sys_tmp459;
	wire        [31:0] w_sys_tmp461;
	wire signed [31:0] w_sys_tmp462;
	wire signed [31:0] w_sys_tmp463;
	wire signed [31:0] w_sys_tmp466;
	wire signed [31:0] w_sys_tmp467;
	wire        [31:0] w_sys_tmp469;
	wire signed [31:0] w_sys_tmp470;
	wire signed [31:0] w_sys_tmp471;
	wire signed [31:0] w_sys_tmp473;
	wire signed [31:0] w_sys_tmp474;
	wire signed [31:0] w_sys_tmp475;
	wire signed [31:0] w_sys_tmp476;
	wire signed [31:0] w_sys_tmp477;
	wire signed [31:0] w_sys_tmp478;
	wire signed [31:0] w_sys_tmp659;
	wire               w_sys_tmp660;
	wire               w_sys_tmp661;
	wire signed [31:0] w_sys_tmp662;
	wire signed [31:0] w_sys_tmp665;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp667;
	wire        [31:0] w_sys_tmp668;
	wire signed [31:0] w_sys_tmp669;
	wire signed [31:0] w_sys_tmp670;
	wire signed [31:0] w_sys_tmp673;
	wire signed [31:0] w_sys_tmp674;
	wire        [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp677;
	wire signed [31:0] w_sys_tmp678;
	wire signed [31:0] w_sys_tmp681;
	wire signed [31:0] w_sys_tmp682;
	wire        [31:0] w_sys_tmp684;
	wire signed [31:0] w_sys_tmp685;
	wire signed [31:0] w_sys_tmp686;
	wire signed [31:0] w_sys_tmp688;
	wire signed [31:0] w_sys_tmp689;
	wire signed [31:0] w_sys_tmp690;
	wire signed [31:0] w_sys_tmp691;
	wire signed [31:0] w_sys_tmp692;
	wire signed [31:0] w_sys_tmp693;
	wire signed [31:0] w_sys_tmp874;
	wire               w_sys_tmp875;
	wire               w_sys_tmp876;
	wire signed [31:0] w_sys_tmp877;
	wire signed [31:0] w_sys_tmp880;
	wire signed [31:0] w_sys_tmp881;
	wire signed [31:0] w_sys_tmp882;
	wire        [31:0] w_sys_tmp883;
	wire signed [31:0] w_sys_tmp884;
	wire signed [31:0] w_sys_tmp885;
	wire signed [31:0] w_sys_tmp888;
	wire signed [31:0] w_sys_tmp889;
	wire        [31:0] w_sys_tmp891;
	wire signed [31:0] w_sys_tmp892;
	wire signed [31:0] w_sys_tmp893;
	wire signed [31:0] w_sys_tmp896;
	wire signed [31:0] w_sys_tmp897;
	wire        [31:0] w_sys_tmp899;
	wire signed [31:0] w_sys_tmp900;
	wire signed [31:0] w_sys_tmp901;
	wire signed [31:0] w_sys_tmp903;
	wire signed [31:0] w_sys_tmp904;
	wire signed [31:0] w_sys_tmp905;
	wire signed [31:0] w_sys_tmp906;
	wire signed [31:0] w_sys_tmp907;
	wire signed [31:0] w_sys_tmp908;
	wire signed [31:0] w_sys_tmp1089;
	wire               w_sys_tmp1090;
	wire               w_sys_tmp1091;
	wire signed [31:0] w_sys_tmp1092;
	wire signed [31:0] w_sys_tmp1093;
	wire               w_sys_tmp1094;
	wire               w_sys_tmp1095;
	wire signed [31:0] w_sys_tmp1096;
	wire signed [31:0] w_sys_tmp1099;
	wire signed [31:0] w_sys_tmp1100;
	wire signed [31:0] w_sys_tmp1101;
	wire        [31:0] w_sys_tmp1102;
	wire signed [31:0] w_sys_tmp1103;
	wire signed [31:0] w_sys_tmp1104;
	wire signed [31:0] w_sys_tmp1107;
	wire signed [31:0] w_sys_tmp1108;
	wire        [31:0] w_sys_tmp1110;
	wire signed [31:0] w_sys_tmp1111;
	wire signed [31:0] w_sys_tmp1112;
	wire signed [31:0] w_sys_tmp1115;
	wire signed [31:0] w_sys_tmp1116;
	wire        [31:0] w_sys_tmp1118;
	wire signed [31:0] w_sys_tmp1119;
	wire signed [31:0] w_sys_tmp1120;
	wire signed [31:0] w_sys_tmp1122;
	wire signed [31:0] w_sys_tmp1123;
	wire signed [31:0] w_sys_tmp1124;
	wire signed [31:0] w_sys_tmp1125;
	wire signed [31:0] w_sys_tmp1126;
	wire signed [31:0] w_sys_tmp1127;
	wire signed [31:0] w_sys_tmp1308;
	wire               w_sys_tmp1309;
	wire               w_sys_tmp1310;
	wire signed [31:0] w_sys_tmp1311;
	wire signed [31:0] w_sys_tmp1314;
	wire signed [31:0] w_sys_tmp1315;
	wire signed [31:0] w_sys_tmp1316;
	wire        [31:0] w_sys_tmp1317;
	wire signed [31:0] w_sys_tmp1318;
	wire signed [31:0] w_sys_tmp1319;
	wire signed [31:0] w_sys_tmp1322;
	wire signed [31:0] w_sys_tmp1323;
	wire        [31:0] w_sys_tmp1325;
	wire signed [31:0] w_sys_tmp1326;
	wire signed [31:0] w_sys_tmp1327;
	wire signed [31:0] w_sys_tmp1330;
	wire signed [31:0] w_sys_tmp1331;
	wire        [31:0] w_sys_tmp1333;
	wire signed [31:0] w_sys_tmp1334;
	wire signed [31:0] w_sys_tmp1335;
	wire signed [31:0] w_sys_tmp1337;
	wire signed [31:0] w_sys_tmp1338;
	wire signed [31:0] w_sys_tmp1339;
	wire signed [31:0] w_sys_tmp1340;
	wire signed [31:0] w_sys_tmp1341;
	wire signed [31:0] w_sys_tmp1342;
	wire signed [31:0] w_sys_tmp1523;
	wire               w_sys_tmp1524;
	wire               w_sys_tmp1525;
	wire signed [31:0] w_sys_tmp1526;
	wire signed [31:0] w_sys_tmp1529;
	wire signed [31:0] w_sys_tmp1530;
	wire signed [31:0] w_sys_tmp1531;
	wire        [31:0] w_sys_tmp1532;
	wire signed [31:0] w_sys_tmp1533;
	wire signed [31:0] w_sys_tmp1534;
	wire signed [31:0] w_sys_tmp1537;
	wire signed [31:0] w_sys_tmp1538;
	wire        [31:0] w_sys_tmp1540;
	wire signed [31:0] w_sys_tmp1541;
	wire signed [31:0] w_sys_tmp1542;
	wire signed [31:0] w_sys_tmp1545;
	wire signed [31:0] w_sys_tmp1546;
	wire        [31:0] w_sys_tmp1548;
	wire signed [31:0] w_sys_tmp1549;
	wire signed [31:0] w_sys_tmp1550;
	wire signed [31:0] w_sys_tmp1552;
	wire signed [31:0] w_sys_tmp1553;
	wire signed [31:0] w_sys_tmp1554;
	wire signed [31:0] w_sys_tmp1555;
	wire signed [31:0] w_sys_tmp1556;
	wire signed [31:0] w_sys_tmp1557;
	wire signed [31:0] w_sys_tmp1738;
	wire               w_sys_tmp1739;
	wire               w_sys_tmp1740;
	wire signed [31:0] w_sys_tmp1741;
	wire signed [31:0] w_sys_tmp1744;
	wire signed [31:0] w_sys_tmp1745;
	wire signed [31:0] w_sys_tmp1746;
	wire        [31:0] w_sys_tmp1747;
	wire signed [31:0] w_sys_tmp1748;
	wire signed [31:0] w_sys_tmp1749;
	wire signed [31:0] w_sys_tmp1752;
	wire signed [31:0] w_sys_tmp1753;
	wire        [31:0] w_sys_tmp1755;
	wire signed [31:0] w_sys_tmp1756;
	wire signed [31:0] w_sys_tmp1757;
	wire signed [31:0] w_sys_tmp1760;
	wire signed [31:0] w_sys_tmp1761;
	wire        [31:0] w_sys_tmp1763;
	wire signed [31:0] w_sys_tmp1764;
	wire signed [31:0] w_sys_tmp1765;
	wire signed [31:0] w_sys_tmp1767;
	wire signed [31:0] w_sys_tmp1768;
	wire signed [31:0] w_sys_tmp1769;
	wire signed [31:0] w_sys_tmp1770;
	wire signed [31:0] w_sys_tmp1771;
	wire signed [31:0] w_sys_tmp1772;
	wire signed [31:0] w_sys_tmp1953;
	wire               w_sys_tmp1954;
	wire               w_sys_tmp1955;
	wire signed [31:0] w_sys_tmp1956;
	wire signed [31:0] w_sys_tmp1957;
	wire               w_sys_tmp1958;
	wire               w_sys_tmp1959;
	wire signed [31:0] w_sys_tmp1960;
	wire signed [31:0] w_sys_tmp1963;
	wire signed [31:0] w_sys_tmp1964;
	wire signed [31:0] w_sys_tmp1965;
	wire        [31:0] w_sys_tmp1966;
	wire signed [31:0] w_sys_tmp1967;
	wire signed [31:0] w_sys_tmp1968;
	wire signed [31:0] w_sys_tmp1971;
	wire signed [31:0] w_sys_tmp1972;
	wire        [31:0] w_sys_tmp1974;
	wire signed [31:0] w_sys_tmp1975;
	wire signed [31:0] w_sys_tmp1976;
	wire signed [31:0] w_sys_tmp1979;
	wire signed [31:0] w_sys_tmp1980;
	wire        [31:0] w_sys_tmp1982;
	wire signed [31:0] w_sys_tmp1983;
	wire signed [31:0] w_sys_tmp1984;
	wire signed [31:0] w_sys_tmp1986;
	wire signed [31:0] w_sys_tmp1987;
	wire signed [31:0] w_sys_tmp1988;
	wire signed [31:0] w_sys_tmp1989;
	wire signed [31:0] w_sys_tmp1990;
	wire signed [31:0] w_sys_tmp1991;
	wire signed [31:0] w_sys_tmp2172;
	wire               w_sys_tmp2173;
	wire               w_sys_tmp2174;
	wire signed [31:0] w_sys_tmp2175;
	wire signed [31:0] w_sys_tmp2178;
	wire signed [31:0] w_sys_tmp2179;
	wire signed [31:0] w_sys_tmp2180;
	wire        [31:0] w_sys_tmp2181;
	wire signed [31:0] w_sys_tmp2182;
	wire signed [31:0] w_sys_tmp2183;
	wire signed [31:0] w_sys_tmp2186;
	wire signed [31:0] w_sys_tmp2187;
	wire        [31:0] w_sys_tmp2189;
	wire signed [31:0] w_sys_tmp2190;
	wire signed [31:0] w_sys_tmp2191;
	wire signed [31:0] w_sys_tmp2194;
	wire signed [31:0] w_sys_tmp2195;
	wire        [31:0] w_sys_tmp2197;
	wire signed [31:0] w_sys_tmp2198;
	wire signed [31:0] w_sys_tmp2199;
	wire signed [31:0] w_sys_tmp2201;
	wire signed [31:0] w_sys_tmp2202;
	wire signed [31:0] w_sys_tmp2203;
	wire signed [31:0] w_sys_tmp2204;
	wire signed [31:0] w_sys_tmp2205;
	wire signed [31:0] w_sys_tmp2206;
	wire signed [31:0] w_sys_tmp2387;
	wire               w_sys_tmp2388;
	wire               w_sys_tmp2389;
	wire signed [31:0] w_sys_tmp2390;
	wire signed [31:0] w_sys_tmp2393;
	wire signed [31:0] w_sys_tmp2394;
	wire signed [31:0] w_sys_tmp2395;
	wire        [31:0] w_sys_tmp2396;
	wire signed [31:0] w_sys_tmp2397;
	wire signed [31:0] w_sys_tmp2398;
	wire signed [31:0] w_sys_tmp2401;
	wire signed [31:0] w_sys_tmp2402;
	wire        [31:0] w_sys_tmp2404;
	wire signed [31:0] w_sys_tmp2405;
	wire signed [31:0] w_sys_tmp2406;
	wire signed [31:0] w_sys_tmp2409;
	wire signed [31:0] w_sys_tmp2410;
	wire        [31:0] w_sys_tmp2412;
	wire signed [31:0] w_sys_tmp2413;
	wire signed [31:0] w_sys_tmp2414;
	wire signed [31:0] w_sys_tmp2416;
	wire signed [31:0] w_sys_tmp2417;
	wire signed [31:0] w_sys_tmp2418;
	wire signed [31:0] w_sys_tmp2419;
	wire signed [31:0] w_sys_tmp2420;
	wire signed [31:0] w_sys_tmp2421;
	wire signed [31:0] w_sys_tmp2602;
	wire               w_sys_tmp2603;
	wire               w_sys_tmp2604;
	wire signed [31:0] w_sys_tmp2605;
	wire signed [31:0] w_sys_tmp2608;
	wire signed [31:0] w_sys_tmp2609;
	wire signed [31:0] w_sys_tmp2610;
	wire        [31:0] w_sys_tmp2611;
	wire signed [31:0] w_sys_tmp2612;
	wire signed [31:0] w_sys_tmp2613;
	wire signed [31:0] w_sys_tmp2616;
	wire signed [31:0] w_sys_tmp2617;
	wire        [31:0] w_sys_tmp2619;
	wire signed [31:0] w_sys_tmp2620;
	wire signed [31:0] w_sys_tmp2621;
	wire signed [31:0] w_sys_tmp2624;
	wire signed [31:0] w_sys_tmp2625;
	wire        [31:0] w_sys_tmp2627;
	wire signed [31:0] w_sys_tmp2628;
	wire signed [31:0] w_sys_tmp2629;
	wire signed [31:0] w_sys_tmp2631;
	wire signed [31:0] w_sys_tmp2632;
	wire signed [31:0] w_sys_tmp2633;
	wire signed [31:0] w_sys_tmp2634;
	wire signed [31:0] w_sys_tmp2635;
	wire signed [31:0] w_sys_tmp2636;
	wire signed [31:0] w_sys_tmp2817;
	wire               w_sys_tmp2818;
	wire               w_sys_tmp2819;
	wire signed [31:0] w_sys_tmp2820;
	wire signed [31:0] w_sys_tmp2821;
	wire               w_sys_tmp2822;
	wire               w_sys_tmp2823;
	wire signed [31:0] w_sys_tmp2824;
	wire signed [31:0] w_sys_tmp2827;
	wire signed [31:0] w_sys_tmp2828;
	wire signed [31:0] w_sys_tmp2829;
	wire        [31:0] w_sys_tmp2830;
	wire signed [31:0] w_sys_tmp2831;
	wire signed [31:0] w_sys_tmp2832;
	wire signed [31:0] w_sys_tmp2835;
	wire signed [31:0] w_sys_tmp2836;
	wire        [31:0] w_sys_tmp2838;
	wire signed [31:0] w_sys_tmp2839;
	wire signed [31:0] w_sys_tmp2840;
	wire signed [31:0] w_sys_tmp2843;
	wire signed [31:0] w_sys_tmp2844;
	wire        [31:0] w_sys_tmp2846;
	wire signed [31:0] w_sys_tmp2847;
	wire signed [31:0] w_sys_tmp2848;
	wire signed [31:0] w_sys_tmp2850;
	wire signed [31:0] w_sys_tmp2851;
	wire signed [31:0] w_sys_tmp2852;
	wire signed [31:0] w_sys_tmp2853;
	wire signed [31:0] w_sys_tmp2854;
	wire signed [31:0] w_sys_tmp2855;
	wire signed [31:0] w_sys_tmp3036;
	wire               w_sys_tmp3037;
	wire               w_sys_tmp3038;
	wire signed [31:0] w_sys_tmp3039;
	wire signed [31:0] w_sys_tmp3042;
	wire signed [31:0] w_sys_tmp3043;
	wire signed [31:0] w_sys_tmp3044;
	wire        [31:0] w_sys_tmp3045;
	wire signed [31:0] w_sys_tmp3046;
	wire signed [31:0] w_sys_tmp3047;
	wire signed [31:0] w_sys_tmp3050;
	wire signed [31:0] w_sys_tmp3051;
	wire        [31:0] w_sys_tmp3053;
	wire signed [31:0] w_sys_tmp3054;
	wire signed [31:0] w_sys_tmp3055;
	wire signed [31:0] w_sys_tmp3058;
	wire signed [31:0] w_sys_tmp3059;
	wire        [31:0] w_sys_tmp3061;
	wire signed [31:0] w_sys_tmp3062;
	wire signed [31:0] w_sys_tmp3063;
	wire signed [31:0] w_sys_tmp3065;
	wire signed [31:0] w_sys_tmp3066;
	wire signed [31:0] w_sys_tmp3067;
	wire signed [31:0] w_sys_tmp3068;
	wire signed [31:0] w_sys_tmp3069;
	wire signed [31:0] w_sys_tmp3070;
	wire signed [31:0] w_sys_tmp3251;
	wire               w_sys_tmp3252;
	wire               w_sys_tmp3253;
	wire signed [31:0] w_sys_tmp3254;
	wire signed [31:0] w_sys_tmp3257;
	wire signed [31:0] w_sys_tmp3258;
	wire signed [31:0] w_sys_tmp3259;
	wire        [31:0] w_sys_tmp3260;
	wire signed [31:0] w_sys_tmp3261;
	wire signed [31:0] w_sys_tmp3262;
	wire signed [31:0] w_sys_tmp3265;
	wire signed [31:0] w_sys_tmp3266;
	wire        [31:0] w_sys_tmp3268;
	wire signed [31:0] w_sys_tmp3269;
	wire signed [31:0] w_sys_tmp3270;
	wire signed [31:0] w_sys_tmp3273;
	wire signed [31:0] w_sys_tmp3274;
	wire        [31:0] w_sys_tmp3276;
	wire signed [31:0] w_sys_tmp3277;
	wire signed [31:0] w_sys_tmp3278;
	wire signed [31:0] w_sys_tmp3280;
	wire signed [31:0] w_sys_tmp3281;
	wire signed [31:0] w_sys_tmp3282;
	wire signed [31:0] w_sys_tmp3283;
	wire signed [31:0] w_sys_tmp3284;
	wire signed [31:0] w_sys_tmp3285;
	wire signed [31:0] w_sys_tmp3466;
	wire               w_sys_tmp3467;
	wire               w_sys_tmp3468;
	wire signed [31:0] w_sys_tmp3469;
	wire signed [31:0] w_sys_tmp3472;
	wire signed [31:0] w_sys_tmp3473;
	wire signed [31:0] w_sys_tmp3474;
	wire        [31:0] w_sys_tmp3475;
	wire signed [31:0] w_sys_tmp3476;
	wire signed [31:0] w_sys_tmp3477;
	wire signed [31:0] w_sys_tmp3480;
	wire signed [31:0] w_sys_tmp3481;
	wire        [31:0] w_sys_tmp3483;
	wire signed [31:0] w_sys_tmp3484;
	wire signed [31:0] w_sys_tmp3485;
	wire signed [31:0] w_sys_tmp3488;
	wire signed [31:0] w_sys_tmp3489;
	wire        [31:0] w_sys_tmp3491;
	wire signed [31:0] w_sys_tmp3492;
	wire signed [31:0] w_sys_tmp3493;
	wire signed [31:0] w_sys_tmp3495;
	wire signed [31:0] w_sys_tmp3496;
	wire signed [31:0] w_sys_tmp3497;
	wire signed [31:0] w_sys_tmp3498;
	wire signed [31:0] w_sys_tmp3499;
	wire signed [31:0] w_sys_tmp3500;
	wire               w_sys_tmp3681;
	wire               w_sys_tmp3682;
	wire signed [31:0] w_sys_tmp3683;
	wire signed [31:0] w_sys_tmp3684;
	wire               w_sys_tmp3685;
	wire               w_sys_tmp3686;
	wire signed [31:0] w_sys_tmp3687;
	wire signed [31:0] w_sys_tmp3690;
	wire signed [31:0] w_sys_tmp3691;
	wire        [31:0] w_sys_tmp3692;
	wire signed [31:0] w_sys_tmp3696;
	wire signed [31:0] w_sys_tmp3697;
	wire        [31:0] w_sys_tmp3698;
	wire signed [31:0] w_sys_tmp3702;
	wire signed [31:0] w_sys_tmp3703;
	wire signed [31:0] w_sys_tmp3707;
	wire signed [31:0] w_sys_tmp3708;
	wire signed [31:0] w_sys_tmp3713;
	wire signed [31:0] w_sys_tmp3714;
	wire signed [31:0] w_sys_tmp3718;
	wire signed [31:0] w_sys_tmp3719;
	wire        [31:0] w_sys_tmp3720;
	wire signed [31:0] w_sys_tmp3723;
	wire signed [31:0] w_sys_tmp3724;
	wire               w_sys_tmp3725;
	wire               w_sys_tmp3726;
	wire signed [31:0] w_sys_tmp3727;
	wire signed [31:0] w_sys_tmp3730;
	wire signed [31:0] w_sys_tmp3731;
	wire        [31:0] w_sys_tmp3732;
	wire signed [31:0] w_sys_tmp3736;
	wire signed [31:0] w_sys_tmp3737;
	wire        [31:0] w_sys_tmp3738;
	wire signed [31:0] w_sys_tmp3742;
	wire signed [31:0] w_sys_tmp3743;
	wire signed [31:0] w_sys_tmp3747;
	wire signed [31:0] w_sys_tmp3748;
	wire signed [31:0] w_sys_tmp3753;
	wire signed [31:0] w_sys_tmp3754;
	wire signed [31:0] w_sys_tmp3758;
	wire signed [31:0] w_sys_tmp3759;
	wire        [31:0] w_sys_tmp3760;
	wire signed [31:0] w_sys_tmp3763;
	wire signed [31:0] w_sys_tmp3764;
	wire               w_sys_tmp3765;
	wire               w_sys_tmp3766;
	wire signed [31:0] w_sys_tmp3767;
	wire signed [31:0] w_sys_tmp3770;
	wire signed [31:0] w_sys_tmp3771;
	wire        [31:0] w_sys_tmp3772;
	wire signed [31:0] w_sys_tmp3776;
	wire signed [31:0] w_sys_tmp3777;
	wire        [31:0] w_sys_tmp3778;
	wire signed [31:0] w_sys_tmp3782;
	wire signed [31:0] w_sys_tmp3783;
	wire signed [31:0] w_sys_tmp3787;
	wire signed [31:0] w_sys_tmp3788;
	wire signed [31:0] w_sys_tmp3793;
	wire signed [31:0] w_sys_tmp3794;
	wire signed [31:0] w_sys_tmp3798;
	wire signed [31:0] w_sys_tmp3799;
	wire        [31:0] w_sys_tmp3800;
	wire signed [31:0] w_sys_tmp3803;
	wire signed [31:0] w_sys_tmp3804;
	wire               w_sys_tmp3805;
	wire               w_sys_tmp3806;
	wire signed [31:0] w_sys_tmp3807;
	wire signed [31:0] w_sys_tmp3810;
	wire signed [31:0] w_sys_tmp3811;
	wire        [31:0] w_sys_tmp3812;
	wire signed [31:0] w_sys_tmp3816;
	wire signed [31:0] w_sys_tmp3817;
	wire        [31:0] w_sys_tmp3818;
	wire signed [31:0] w_sys_tmp3822;
	wire signed [31:0] w_sys_tmp3823;
	wire signed [31:0] w_sys_tmp3827;
	wire signed [31:0] w_sys_tmp3828;
	wire signed [31:0] w_sys_tmp3833;
	wire signed [31:0] w_sys_tmp3834;
	wire signed [31:0] w_sys_tmp3838;
	wire signed [31:0] w_sys_tmp3839;
	wire        [31:0] w_sys_tmp3840;
	wire signed [31:0] w_sys_tmp3843;
	wire signed [31:0] w_sys_tmp3844;
	wire               w_sys_tmp3845;
	wire               w_sys_tmp3846;
	wire signed [31:0] w_sys_tmp3847;
	wire signed [31:0] w_sys_tmp3850;
	wire signed [31:0] w_sys_tmp3851;
	wire signed [31:0] w_sys_tmp3852;
	wire signed [31:0] w_sys_tmp3853;
	wire        [31:0] w_sys_tmp3854;
	wire signed [31:0] w_sys_tmp3855;
	wire signed [31:0] w_sys_tmp3856;
	wire signed [31:0] w_sys_tmp3860;
	wire signed [31:0] w_sys_tmp3861;
	wire signed [31:0] w_sys_tmp3863;
	wire        [31:0] w_sys_tmp3864;
	wire signed [31:0] w_sys_tmp3865;
	wire signed [31:0] w_sys_tmp3866;
	wire signed [31:0] w_sys_tmp3870;
	wire signed [31:0] w_sys_tmp3871;
	wire signed [31:0] w_sys_tmp3873;
	wire signed [31:0] w_sys_tmp3874;
	wire signed [31:0] w_sys_tmp3875;
	wire signed [31:0] w_sys_tmp3879;
	wire signed [31:0] w_sys_tmp3880;
	wire signed [31:0] w_sys_tmp3882;
	wire signed [31:0] w_sys_tmp3884;
	wire signed [31:0] w_sys_tmp3885;
	wire signed [31:0] w_sys_tmp3889;
	wire signed [31:0] w_sys_tmp3890;
	wire signed [31:0] w_sys_tmp3892;
	wire signed [31:0] w_sys_tmp3893;
	wire signed [31:0] w_sys_tmp3894;
	wire signed [31:0] w_sys_tmp3898;
	wire signed [31:0] w_sys_tmp3899;
	wire signed [31:0] w_sys_tmp3901;
	wire        [31:0] w_sys_tmp3902;
	wire signed [31:0] w_sys_tmp3903;
	wire signed [31:0] w_sys_tmp3904;
	wire signed [31:0] w_sys_tmp3907;
	wire signed [31:0] w_sys_tmp3908;
	wire signed [31:0] w_sys_tmp3909;
	wire signed [31:0] w_sys_tmp3910;
	wire signed [31:0] w_sys_tmp3911;
	wire signed [31:0] w_sys_tmp3912;
	wire signed [31:0] w_sys_tmp3913;
	wire signed [31:0] w_sys_tmp3914;
	wire signed [31:0] w_sys_tmp3915;
	wire signed [31:0] w_sys_tmp3916;
	wire signed [31:0] w_sys_tmp3917;
	wire signed [31:0] w_sys_tmp3918;
	wire signed [31:0] w_sys_tmp4345;
	wire               w_sys_tmp4346;
	wire               w_sys_tmp4347;
	wire signed [31:0] w_sys_tmp4348;
	wire signed [31:0] w_sys_tmp4351;
	wire signed [31:0] w_sys_tmp4352;
	wire signed [31:0] w_sys_tmp4353;
	wire signed [31:0] w_sys_tmp4354;
	wire        [31:0] w_sys_tmp4355;
	wire signed [31:0] w_sys_tmp4356;
	wire signed [31:0] w_sys_tmp4357;
	wire signed [31:0] w_sys_tmp4361;
	wire signed [31:0] w_sys_tmp4362;
	wire signed [31:0] w_sys_tmp4364;
	wire        [31:0] w_sys_tmp4365;
	wire signed [31:0] w_sys_tmp4366;
	wire signed [31:0] w_sys_tmp4367;
	wire signed [31:0] w_sys_tmp4371;
	wire signed [31:0] w_sys_tmp4372;
	wire signed [31:0] w_sys_tmp4374;
	wire signed [31:0] w_sys_tmp4375;
	wire signed [31:0] w_sys_tmp4376;
	wire signed [31:0] w_sys_tmp4380;
	wire signed [31:0] w_sys_tmp4381;
	wire signed [31:0] w_sys_tmp4383;
	wire signed [31:0] w_sys_tmp4385;
	wire signed [31:0] w_sys_tmp4386;
	wire signed [31:0] w_sys_tmp4390;
	wire signed [31:0] w_sys_tmp4391;
	wire signed [31:0] w_sys_tmp4393;
	wire signed [31:0] w_sys_tmp4394;
	wire signed [31:0] w_sys_tmp4395;
	wire signed [31:0] w_sys_tmp4399;
	wire signed [31:0] w_sys_tmp4400;
	wire signed [31:0] w_sys_tmp4402;
	wire        [31:0] w_sys_tmp4403;
	wire signed [31:0] w_sys_tmp4404;
	wire signed [31:0] w_sys_tmp4405;
	wire signed [31:0] w_sys_tmp4408;
	wire signed [31:0] w_sys_tmp4409;
	wire signed [31:0] w_sys_tmp4410;
	wire signed [31:0] w_sys_tmp4411;
	wire signed [31:0] w_sys_tmp4412;
	wire signed [31:0] w_sys_tmp4413;
	wire signed [31:0] w_sys_tmp4414;
	wire signed [31:0] w_sys_tmp4415;
	wire signed [31:0] w_sys_tmp4416;
	wire signed [31:0] w_sys_tmp4417;
	wire signed [31:0] w_sys_tmp4418;
	wire signed [31:0] w_sys_tmp4419;
	wire signed [31:0] w_sys_tmp4846;
	wire               w_sys_tmp4847;
	wire               w_sys_tmp4848;
	wire signed [31:0] w_sys_tmp4849;
	wire signed [31:0] w_sys_tmp4852;
	wire signed [31:0] w_sys_tmp4853;
	wire signed [31:0] w_sys_tmp4854;
	wire signed [31:0] w_sys_tmp4855;
	wire        [31:0] w_sys_tmp4856;
	wire signed [31:0] w_sys_tmp4857;
	wire signed [31:0] w_sys_tmp4858;
	wire signed [31:0] w_sys_tmp4862;
	wire signed [31:0] w_sys_tmp4863;
	wire signed [31:0] w_sys_tmp4865;
	wire        [31:0] w_sys_tmp4866;
	wire signed [31:0] w_sys_tmp4867;
	wire signed [31:0] w_sys_tmp4868;
	wire signed [31:0] w_sys_tmp4872;
	wire signed [31:0] w_sys_tmp4873;
	wire signed [31:0] w_sys_tmp4875;
	wire signed [31:0] w_sys_tmp4876;
	wire signed [31:0] w_sys_tmp4877;
	wire signed [31:0] w_sys_tmp4881;
	wire signed [31:0] w_sys_tmp4882;
	wire signed [31:0] w_sys_tmp4884;
	wire signed [31:0] w_sys_tmp4886;
	wire signed [31:0] w_sys_tmp4887;
	wire signed [31:0] w_sys_tmp4891;
	wire signed [31:0] w_sys_tmp4892;
	wire signed [31:0] w_sys_tmp4894;
	wire signed [31:0] w_sys_tmp4895;
	wire signed [31:0] w_sys_tmp4896;
	wire signed [31:0] w_sys_tmp4900;
	wire signed [31:0] w_sys_tmp4901;
	wire signed [31:0] w_sys_tmp4903;
	wire        [31:0] w_sys_tmp4904;
	wire signed [31:0] w_sys_tmp4905;
	wire signed [31:0] w_sys_tmp4906;
	wire signed [31:0] w_sys_tmp4909;
	wire signed [31:0] w_sys_tmp4910;
	wire signed [31:0] w_sys_tmp4911;
	wire signed [31:0] w_sys_tmp4912;
	wire signed [31:0] w_sys_tmp4913;
	wire signed [31:0] w_sys_tmp4914;
	wire signed [31:0] w_sys_tmp4915;
	wire signed [31:0] w_sys_tmp4916;
	wire signed [31:0] w_sys_tmp4917;
	wire signed [31:0] w_sys_tmp4918;
	wire signed [31:0] w_sys_tmp4919;
	wire signed [31:0] w_sys_tmp4920;
	wire signed [31:0] w_sys_tmp5347;
	wire               w_sys_tmp5348;
	wire               w_sys_tmp5349;
	wire signed [31:0] w_sys_tmp5350;
	wire signed [31:0] w_sys_tmp5353;
	wire signed [31:0] w_sys_tmp5354;
	wire signed [31:0] w_sys_tmp5355;
	wire signed [31:0] w_sys_tmp5356;
	wire        [31:0] w_sys_tmp5357;
	wire signed [31:0] w_sys_tmp5358;
	wire signed [31:0] w_sys_tmp5359;
	wire signed [31:0] w_sys_tmp5363;
	wire signed [31:0] w_sys_tmp5364;
	wire signed [31:0] w_sys_tmp5366;
	wire        [31:0] w_sys_tmp5367;
	wire signed [31:0] w_sys_tmp5368;
	wire signed [31:0] w_sys_tmp5369;
	wire signed [31:0] w_sys_tmp5373;
	wire signed [31:0] w_sys_tmp5374;
	wire signed [31:0] w_sys_tmp5376;
	wire signed [31:0] w_sys_tmp5377;
	wire signed [31:0] w_sys_tmp5378;
	wire signed [31:0] w_sys_tmp5382;
	wire signed [31:0] w_sys_tmp5383;
	wire signed [31:0] w_sys_tmp5385;
	wire signed [31:0] w_sys_tmp5387;
	wire signed [31:0] w_sys_tmp5388;
	wire signed [31:0] w_sys_tmp5392;
	wire signed [31:0] w_sys_tmp5393;
	wire signed [31:0] w_sys_tmp5395;
	wire signed [31:0] w_sys_tmp5396;
	wire signed [31:0] w_sys_tmp5397;
	wire signed [31:0] w_sys_tmp5401;
	wire signed [31:0] w_sys_tmp5402;
	wire signed [31:0] w_sys_tmp5404;
	wire        [31:0] w_sys_tmp5405;
	wire signed [31:0] w_sys_tmp5406;
	wire signed [31:0] w_sys_tmp5407;
	wire signed [31:0] w_sys_tmp5410;
	wire signed [31:0] w_sys_tmp5411;
	wire signed [31:0] w_sys_tmp5412;
	wire signed [31:0] w_sys_tmp5413;
	wire signed [31:0] w_sys_tmp5414;
	wire signed [31:0] w_sys_tmp5415;
	wire signed [31:0] w_sys_tmp5416;
	wire signed [31:0] w_sys_tmp5417;
	wire signed [31:0] w_sys_tmp5418;
	wire signed [31:0] w_sys_tmp5419;
	wire signed [31:0] w_sys_tmp5420;
	wire signed [31:0] w_sys_tmp5421;
	wire signed [31:0] w_sys_tmp5848;
	wire               w_sys_tmp5849;
	wire               w_sys_tmp5850;
	wire signed [31:0] w_sys_tmp5851;
	wire signed [31:0] w_sys_tmp5852;
	wire signed [31:0] w_sys_tmp5853;
	wire               w_sys_tmp5854;
	wire               w_sys_tmp5855;
	wire signed [31:0] w_sys_tmp5856;
	wire signed [31:0] w_sys_tmp5859;
	wire signed [31:0] w_sys_tmp5860;
	wire signed [31:0] w_sys_tmp5861;
	wire        [31:0] w_sys_tmp5862;
	wire signed [31:0] w_sys_tmp5863;
	wire signed [31:0] w_sys_tmp5864;
	wire signed [31:0] w_sys_tmp5866;
	wire signed [31:0] w_sys_tmp5867;
	wire signed [31:0] w_sys_tmp5928;
	wire               w_sys_tmp5929;
	wire               w_sys_tmp5930;
	wire signed [31:0] w_sys_tmp5931;
	wire signed [31:0] w_sys_tmp5934;
	wire signed [31:0] w_sys_tmp5935;
	wire signed [31:0] w_sys_tmp5936;
	wire        [31:0] w_sys_tmp5937;
	wire signed [31:0] w_sys_tmp5938;
	wire signed [31:0] w_sys_tmp5939;
	wire signed [31:0] w_sys_tmp5941;
	wire signed [31:0] w_sys_tmp5942;
	wire signed [31:0] w_sys_tmp6003;
	wire               w_sys_tmp6004;
	wire               w_sys_tmp6005;
	wire signed [31:0] w_sys_tmp6006;
	wire signed [31:0] w_sys_tmp6009;
	wire signed [31:0] w_sys_tmp6010;
	wire signed [31:0] w_sys_tmp6011;
	wire        [31:0] w_sys_tmp6012;
	wire signed [31:0] w_sys_tmp6013;
	wire signed [31:0] w_sys_tmp6014;
	wire signed [31:0] w_sys_tmp6016;
	wire signed [31:0] w_sys_tmp6017;
	wire signed [31:0] w_sys_tmp6078;
	wire               w_sys_tmp6079;
	wire               w_sys_tmp6080;
	wire signed [31:0] w_sys_tmp6081;
	wire signed [31:0] w_sys_tmp6084;
	wire signed [31:0] w_sys_tmp6085;
	wire signed [31:0] w_sys_tmp6086;
	wire        [31:0] w_sys_tmp6087;
	wire signed [31:0] w_sys_tmp6088;
	wire signed [31:0] w_sys_tmp6089;
	wire signed [31:0] w_sys_tmp6091;
	wire signed [31:0] w_sys_tmp6092;
	wire signed [31:0] w_sys_tmp6153;
	wire               w_sys_tmp6154;
	wire               w_sys_tmp6155;
	wire signed [31:0] w_sys_tmp6156;
	wire signed [31:0] w_sys_tmp6157;
	wire signed [31:0] w_sys_tmp6158;
	wire               w_sys_tmp6159;
	wire               w_sys_tmp6160;
	wire signed [31:0] w_sys_tmp6161;
	wire signed [31:0] w_sys_tmp6164;
	wire signed [31:0] w_sys_tmp6165;
	wire signed [31:0] w_sys_tmp6166;
	wire        [31:0] w_sys_tmp6167;
	wire signed [31:0] w_sys_tmp6168;
	wire signed [31:0] w_sys_tmp6169;
	wire signed [31:0] w_sys_tmp6171;
	wire signed [31:0] w_sys_tmp6172;
	wire signed [31:0] w_sys_tmp6233;
	wire               w_sys_tmp6234;
	wire               w_sys_tmp6235;
	wire signed [31:0] w_sys_tmp6236;
	wire signed [31:0] w_sys_tmp6239;
	wire signed [31:0] w_sys_tmp6240;
	wire signed [31:0] w_sys_tmp6241;
	wire        [31:0] w_sys_tmp6242;
	wire signed [31:0] w_sys_tmp6243;
	wire signed [31:0] w_sys_tmp6244;
	wire signed [31:0] w_sys_tmp6246;
	wire signed [31:0] w_sys_tmp6247;
	wire signed [31:0] w_sys_tmp6308;
	wire               w_sys_tmp6309;
	wire               w_sys_tmp6310;
	wire signed [31:0] w_sys_tmp6311;
	wire signed [31:0] w_sys_tmp6314;
	wire signed [31:0] w_sys_tmp6315;
	wire signed [31:0] w_sys_tmp6316;
	wire        [31:0] w_sys_tmp6317;
	wire signed [31:0] w_sys_tmp6318;
	wire signed [31:0] w_sys_tmp6319;
	wire signed [31:0] w_sys_tmp6321;
	wire signed [31:0] w_sys_tmp6322;
	wire signed [31:0] w_sys_tmp6383;
	wire               w_sys_tmp6384;
	wire               w_sys_tmp6385;
	wire signed [31:0] w_sys_tmp6386;
	wire signed [31:0] w_sys_tmp6389;
	wire signed [31:0] w_sys_tmp6390;
	wire signed [31:0] w_sys_tmp6391;
	wire        [31:0] w_sys_tmp6392;
	wire signed [31:0] w_sys_tmp6393;
	wire signed [31:0] w_sys_tmp6394;
	wire signed [31:0] w_sys_tmp6396;
	wire signed [31:0] w_sys_tmp6397;
	wire signed [31:0] w_sys_tmp6458;
	wire               w_sys_tmp6459;
	wire               w_sys_tmp6460;
	wire signed [31:0] w_sys_tmp6461;
	wire signed [31:0] w_sys_tmp6462;
	wire signed [31:0] w_sys_tmp6463;
	wire               w_sys_tmp6464;
	wire               w_sys_tmp6465;
	wire signed [31:0] w_sys_tmp6466;
	wire signed [31:0] w_sys_tmp6469;
	wire signed [31:0] w_sys_tmp6470;
	wire signed [31:0] w_sys_tmp6471;
	wire        [31:0] w_sys_tmp6472;
	wire signed [31:0] w_sys_tmp6473;
	wire signed [31:0] w_sys_tmp6474;
	wire signed [31:0] w_sys_tmp6476;
	wire signed [31:0] w_sys_tmp6477;
	wire signed [31:0] w_sys_tmp6538;
	wire               w_sys_tmp6539;
	wire               w_sys_tmp6540;
	wire signed [31:0] w_sys_tmp6541;
	wire signed [31:0] w_sys_tmp6544;
	wire signed [31:0] w_sys_tmp6545;
	wire signed [31:0] w_sys_tmp6546;
	wire        [31:0] w_sys_tmp6547;
	wire signed [31:0] w_sys_tmp6548;
	wire signed [31:0] w_sys_tmp6549;
	wire signed [31:0] w_sys_tmp6551;
	wire signed [31:0] w_sys_tmp6552;
	wire signed [31:0] w_sys_tmp6613;
	wire               w_sys_tmp6614;
	wire               w_sys_tmp6615;
	wire signed [31:0] w_sys_tmp6616;
	wire signed [31:0] w_sys_tmp6619;
	wire signed [31:0] w_sys_tmp6620;
	wire signed [31:0] w_sys_tmp6621;
	wire        [31:0] w_sys_tmp6622;
	wire signed [31:0] w_sys_tmp6623;
	wire signed [31:0] w_sys_tmp6624;
	wire signed [31:0] w_sys_tmp6626;
	wire signed [31:0] w_sys_tmp6627;
	wire signed [31:0] w_sys_tmp6688;
	wire               w_sys_tmp6689;
	wire               w_sys_tmp6690;
	wire signed [31:0] w_sys_tmp6691;
	wire signed [31:0] w_sys_tmp6694;
	wire signed [31:0] w_sys_tmp6695;
	wire signed [31:0] w_sys_tmp6696;
	wire        [31:0] w_sys_tmp6697;
	wire signed [31:0] w_sys_tmp6698;
	wire signed [31:0] w_sys_tmp6699;
	wire signed [31:0] w_sys_tmp6701;
	wire signed [31:0] w_sys_tmp6702;
	wire signed [31:0] w_sys_tmp6763;
	wire               w_sys_tmp6764;
	wire               w_sys_tmp6765;
	wire signed [31:0] w_sys_tmp6766;
	wire signed [31:0] w_sys_tmp6767;
	wire signed [31:0] w_sys_tmp6768;
	wire               w_sys_tmp6769;
	wire               w_sys_tmp6770;
	wire signed [31:0] w_sys_tmp6771;
	wire signed [31:0] w_sys_tmp6774;
	wire signed [31:0] w_sys_tmp6775;
	wire signed [31:0] w_sys_tmp6776;
	wire        [31:0] w_sys_tmp6777;
	wire signed [31:0] w_sys_tmp6778;
	wire signed [31:0] w_sys_tmp6779;
	wire signed [31:0] w_sys_tmp6781;
	wire signed [31:0] w_sys_tmp6782;
	wire signed [31:0] w_sys_tmp6843;
	wire               w_sys_tmp6844;
	wire               w_sys_tmp6845;
	wire signed [31:0] w_sys_tmp6846;
	wire signed [31:0] w_sys_tmp6849;
	wire signed [31:0] w_sys_tmp6850;
	wire signed [31:0] w_sys_tmp6851;
	wire        [31:0] w_sys_tmp6852;
	wire signed [31:0] w_sys_tmp6853;
	wire signed [31:0] w_sys_tmp6854;
	wire signed [31:0] w_sys_tmp6856;
	wire signed [31:0] w_sys_tmp6857;
	wire signed [31:0] w_sys_tmp6918;
	wire               w_sys_tmp6919;
	wire               w_sys_tmp6920;
	wire signed [31:0] w_sys_tmp6921;
	wire signed [31:0] w_sys_tmp6924;
	wire signed [31:0] w_sys_tmp6925;
	wire signed [31:0] w_sys_tmp6926;
	wire        [31:0] w_sys_tmp6927;
	wire signed [31:0] w_sys_tmp6928;
	wire signed [31:0] w_sys_tmp6929;
	wire signed [31:0] w_sys_tmp6931;
	wire signed [31:0] w_sys_tmp6932;
	wire signed [31:0] w_sys_tmp6993;
	wire               w_sys_tmp6994;
	wire               w_sys_tmp6995;
	wire signed [31:0] w_sys_tmp6996;
	wire signed [31:0] w_sys_tmp6999;
	wire signed [31:0] w_sys_tmp7000;
	wire signed [31:0] w_sys_tmp7001;
	wire        [31:0] w_sys_tmp7002;
	wire signed [31:0] w_sys_tmp7003;
	wire signed [31:0] w_sys_tmp7004;
	wire signed [31:0] w_sys_tmp7006;
	wire signed [31:0] w_sys_tmp7007;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 6'h1);
	assign w_fld_T_0_addr_0 = 15'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 15'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 15'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_fld_V_3_addr_0 = 15'sh0;
	assign w_fld_V_3_datain_0 = 32'h0;
	assign w_fld_V_3_r_w_0 = 1'h0;
	assign w_fld_V_3_ce_0 = w_sys_ce;
	assign w_fld_V_3_ce_1 = w_sys_ce;
	assign w_sub09_T_addr = ( (|r_sys_processing_methodID) ? r_sub09_T_addr : 15'sh0 ) ;
	assign w_sub09_T_datain = ( (|r_sys_processing_methodID) ? r_sub09_T_datain : 32'h0 ) ;
	assign w_sub09_T_r_w = ( (|r_sys_processing_methodID) ? r_sub09_T_r_w : 1'h0 ) ;
	assign w_sub09_V_addr = ( (|r_sys_processing_methodID) ? r_sub09_V_addr : 15'sh0 ) ;
	assign w_sub09_V_datain = ( (|r_sys_processing_methodID) ? r_sub09_V_datain : 32'h0 ) ;
	assign w_sub09_V_r_w = ( (|r_sys_processing_methodID) ? r_sub09_V_r_w : 1'h0 ) ;
	assign w_sub09_U_addr = ( (|r_sys_processing_methodID) ? r_sub09_U_addr : 15'sh0 ) ;
	assign w_sub09_U_datain = ( (|r_sys_processing_methodID) ? r_sub09_U_datain : 32'h0 ) ;
	assign w_sub09_U_r_w = ( (|r_sys_processing_methodID) ? r_sub09_U_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 15'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_T_addr = ( (|r_sys_processing_methodID) ? r_sub08_T_addr : 15'sh0 ) ;
	assign w_sub08_T_datain = ( (|r_sys_processing_methodID) ? r_sub08_T_datain : 32'h0 ) ;
	assign w_sub08_T_r_w = ( (|r_sys_processing_methodID) ? r_sub08_T_r_w : 1'h0 ) ;
	assign w_sub08_V_addr = ( (|r_sys_processing_methodID) ? r_sub08_V_addr : 15'sh0 ) ;
	assign w_sub08_V_datain = ( (|r_sys_processing_methodID) ? r_sub08_V_datain : 32'h0 ) ;
	assign w_sub08_V_r_w = ( (|r_sys_processing_methodID) ? r_sub08_V_r_w : 1'h0 ) ;
	assign w_sub08_U_addr = ( (|r_sys_processing_methodID) ? r_sub08_U_addr : 15'sh0 ) ;
	assign w_sub08_U_datain = ( (|r_sys_processing_methodID) ? r_sub08_U_datain : 32'h0 ) ;
	assign w_sub08_U_r_w = ( (|r_sys_processing_methodID) ? r_sub08_U_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 15'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub12_T_addr = ( (|r_sys_processing_methodID) ? r_sub12_T_addr : 15'sh0 ) ;
	assign w_sub12_T_datain = ( (|r_sys_processing_methodID) ? r_sub12_T_datain : 32'h0 ) ;
	assign w_sub12_T_r_w = ( (|r_sys_processing_methodID) ? r_sub12_T_r_w : 1'h0 ) ;
	assign w_sub12_V_addr = ( (|r_sys_processing_methodID) ? r_sub12_V_addr : 15'sh0 ) ;
	assign w_sub12_V_datain = ( (|r_sys_processing_methodID) ? r_sub12_V_datain : 32'h0 ) ;
	assign w_sub12_V_r_w = ( (|r_sys_processing_methodID) ? r_sub12_V_r_w : 1'h0 ) ;
	assign w_sub12_U_addr = ( (|r_sys_processing_methodID) ? r_sub12_U_addr : 15'sh0 ) ;
	assign w_sub12_U_datain = ( (|r_sys_processing_methodID) ? r_sub12_U_datain : 32'h0 ) ;
	assign w_sub12_U_r_w = ( (|r_sys_processing_methodID) ? r_sub12_U_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 15'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_T_addr = ( (|r_sys_processing_methodID) ? r_sub03_T_addr : 15'sh0 ) ;
	assign w_sub03_T_datain = ( (|r_sys_processing_methodID) ? r_sub03_T_datain : 32'h0 ) ;
	assign w_sub03_T_r_w = ( (|r_sys_processing_methodID) ? r_sub03_T_r_w : 1'h0 ) ;
	assign w_sub03_V_addr = ( (|r_sys_processing_methodID) ? r_sub03_V_addr : 15'sh0 ) ;
	assign w_sub03_V_datain = ( (|r_sys_processing_methodID) ? r_sub03_V_datain : 32'h0 ) ;
	assign w_sub03_V_r_w = ( (|r_sys_processing_methodID) ? r_sub03_V_r_w : 1'h0 ) ;
	assign w_sub03_U_addr = ( (|r_sys_processing_methodID) ? r_sub03_U_addr : 15'sh0 ) ;
	assign w_sub03_U_datain = ( (|r_sys_processing_methodID) ? r_sub03_U_datain : 32'h0 ) ;
	assign w_sub03_U_r_w = ( (|r_sys_processing_methodID) ? r_sub03_U_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 15'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_T_addr = ( (|r_sys_processing_methodID) ? r_sub02_T_addr : 15'sh0 ) ;
	assign w_sub02_T_datain = ( (|r_sys_processing_methodID) ? r_sub02_T_datain : 32'h0 ) ;
	assign w_sub02_T_r_w = ( (|r_sys_processing_methodID) ? r_sub02_T_r_w : 1'h0 ) ;
	assign w_sub02_V_addr = ( (|r_sys_processing_methodID) ? r_sub02_V_addr : 15'sh0 ) ;
	assign w_sub02_V_datain = ( (|r_sys_processing_methodID) ? r_sub02_V_datain : 32'h0 ) ;
	assign w_sub02_V_r_w = ( (|r_sys_processing_methodID) ? r_sub02_V_r_w : 1'h0 ) ;
	assign w_sub02_U_addr = ( (|r_sys_processing_methodID) ? r_sub02_U_addr : 15'sh0 ) ;
	assign w_sub02_U_datain = ( (|r_sys_processing_methodID) ? r_sub02_U_datain : 32'h0 ) ;
	assign w_sub02_U_r_w = ( (|r_sys_processing_methodID) ? r_sub02_U_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 15'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_T_addr = ( (|r_sys_processing_methodID) ? r_sub11_T_addr : 15'sh0 ) ;
	assign w_sub11_T_datain = ( (|r_sys_processing_methodID) ? r_sub11_T_datain : 32'h0 ) ;
	assign w_sub11_T_r_w = ( (|r_sys_processing_methodID) ? r_sub11_T_r_w : 1'h0 ) ;
	assign w_sub11_V_addr = ( (|r_sys_processing_methodID) ? r_sub11_V_addr : 15'sh0 ) ;
	assign w_sub11_V_datain = ( (|r_sys_processing_methodID) ? r_sub11_V_datain : 32'h0 ) ;
	assign w_sub11_V_r_w = ( (|r_sys_processing_methodID) ? r_sub11_V_r_w : 1'h0 ) ;
	assign w_sub11_U_addr = ( (|r_sys_processing_methodID) ? r_sub11_U_addr : 15'sh0 ) ;
	assign w_sub11_U_datain = ( (|r_sys_processing_methodID) ? r_sub11_U_datain : 32'h0 ) ;
	assign w_sub11_U_r_w = ( (|r_sys_processing_methodID) ? r_sub11_U_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 15'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_T_addr = ( (|r_sys_processing_methodID) ? r_sub14_T_addr : 15'sh0 ) ;
	assign w_sub14_T_datain = ( (|r_sys_processing_methodID) ? r_sub14_T_datain : 32'h0 ) ;
	assign w_sub14_T_r_w = ( (|r_sys_processing_methodID) ? r_sub14_T_r_w : 1'h0 ) ;
	assign w_sub14_V_addr = ( (|r_sys_processing_methodID) ? r_sub14_V_addr : 15'sh0 ) ;
	assign w_sub14_V_datain = ( (|r_sys_processing_methodID) ? r_sub14_V_datain : 32'h0 ) ;
	assign w_sub14_V_r_w = ( (|r_sys_processing_methodID) ? r_sub14_V_r_w : 1'h0 ) ;
	assign w_sub14_U_addr = ( (|r_sys_processing_methodID) ? r_sub14_U_addr : 15'sh0 ) ;
	assign w_sub14_U_datain = ( (|r_sys_processing_methodID) ? r_sub14_U_datain : 32'h0 ) ;
	assign w_sub14_U_r_w = ( (|r_sys_processing_methodID) ? r_sub14_U_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 15'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_T_addr = ( (|r_sys_processing_methodID) ? r_sub01_T_addr : 15'sh0 ) ;
	assign w_sub01_T_datain = ( (|r_sys_processing_methodID) ? r_sub01_T_datain : 32'h0 ) ;
	assign w_sub01_T_r_w = ( (|r_sys_processing_methodID) ? r_sub01_T_r_w : 1'h0 ) ;
	assign w_sub01_V_addr = ( (|r_sys_processing_methodID) ? r_sub01_V_addr : 15'sh0 ) ;
	assign w_sub01_V_datain = ( (|r_sys_processing_methodID) ? r_sub01_V_datain : 32'h0 ) ;
	assign w_sub01_V_r_w = ( (|r_sys_processing_methodID) ? r_sub01_V_r_w : 1'h0 ) ;
	assign w_sub01_U_addr = ( (|r_sys_processing_methodID) ? r_sub01_U_addr : 15'sh0 ) ;
	assign w_sub01_U_datain = ( (|r_sys_processing_methodID) ? r_sub01_U_datain : 32'h0 ) ;
	assign w_sub01_U_r_w = ( (|r_sys_processing_methodID) ? r_sub01_U_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 15'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub13_T_addr = ( (|r_sys_processing_methodID) ? r_sub13_T_addr : 15'sh0 ) ;
	assign w_sub13_T_datain = ( (|r_sys_processing_methodID) ? r_sub13_T_datain : 32'h0 ) ;
	assign w_sub13_T_r_w = ( (|r_sys_processing_methodID) ? r_sub13_T_r_w : 1'h0 ) ;
	assign w_sub13_V_addr = ( (|r_sys_processing_methodID) ? r_sub13_V_addr : 15'sh0 ) ;
	assign w_sub13_V_datain = ( (|r_sys_processing_methodID) ? r_sub13_V_datain : 32'h0 ) ;
	assign w_sub13_V_r_w = ( (|r_sys_processing_methodID) ? r_sub13_V_r_w : 1'h0 ) ;
	assign w_sub13_U_addr = ( (|r_sys_processing_methodID) ? r_sub13_U_addr : 15'sh0 ) ;
	assign w_sub13_U_datain = ( (|r_sys_processing_methodID) ? r_sub13_U_datain : 32'h0 ) ;
	assign w_sub13_U_r_w = ( (|r_sys_processing_methodID) ? r_sub13_U_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 15'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub00_T_addr = ( (|r_sys_processing_methodID) ? r_sub00_T_addr : 15'sh0 ) ;
	assign w_sub00_T_datain = ( (|r_sys_processing_methodID) ? r_sub00_T_datain : 32'h0 ) ;
	assign w_sub00_T_r_w = ( (|r_sys_processing_methodID) ? r_sub00_T_r_w : 1'h0 ) ;
	assign w_sub00_V_addr = ( (|r_sys_processing_methodID) ? r_sub00_V_addr : 15'sh0 ) ;
	assign w_sub00_V_datain = ( (|r_sys_processing_methodID) ? r_sub00_V_datain : 32'h0 ) ;
	assign w_sub00_V_r_w = ( (|r_sys_processing_methodID) ? r_sub00_V_r_w : 1'h0 ) ;
	assign w_sub00_U_addr = ( (|r_sys_processing_methodID) ? r_sub00_U_addr : 15'sh0 ) ;
	assign w_sub00_U_datain = ( (|r_sys_processing_methodID) ? r_sub00_U_datain : 32'h0 ) ;
	assign w_sub00_U_r_w = ( (|r_sys_processing_methodID) ? r_sub00_U_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 15'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_T_addr = ( (|r_sys_processing_methodID) ? r_sub07_T_addr : 15'sh0 ) ;
	assign w_sub07_T_datain = ( (|r_sys_processing_methodID) ? r_sub07_T_datain : 32'h0 ) ;
	assign w_sub07_T_r_w = ( (|r_sys_processing_methodID) ? r_sub07_T_r_w : 1'h0 ) ;
	assign w_sub07_V_addr = ( (|r_sys_processing_methodID) ? r_sub07_V_addr : 15'sh0 ) ;
	assign w_sub07_V_datain = ( (|r_sys_processing_methodID) ? r_sub07_V_datain : 32'h0 ) ;
	assign w_sub07_V_r_w = ( (|r_sys_processing_methodID) ? r_sub07_V_r_w : 1'h0 ) ;
	assign w_sub07_U_addr = ( (|r_sys_processing_methodID) ? r_sub07_U_addr : 15'sh0 ) ;
	assign w_sub07_U_datain = ( (|r_sys_processing_methodID) ? r_sub07_U_datain : 32'h0 ) ;
	assign w_sub07_U_r_w = ( (|r_sys_processing_methodID) ? r_sub07_U_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 15'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_T_addr = ( (|r_sys_processing_methodID) ? r_sub06_T_addr : 15'sh0 ) ;
	assign w_sub06_T_datain = ( (|r_sys_processing_methodID) ? r_sub06_T_datain : 32'h0 ) ;
	assign w_sub06_T_r_w = ( (|r_sys_processing_methodID) ? r_sub06_T_r_w : 1'h0 ) ;
	assign w_sub06_V_addr = ( (|r_sys_processing_methodID) ? r_sub06_V_addr : 15'sh0 ) ;
	assign w_sub06_V_datain = ( (|r_sys_processing_methodID) ? r_sub06_V_datain : 32'h0 ) ;
	assign w_sub06_V_r_w = ( (|r_sys_processing_methodID) ? r_sub06_V_r_w : 1'h0 ) ;
	assign w_sub06_U_addr = ( (|r_sys_processing_methodID) ? r_sub06_U_addr : 15'sh0 ) ;
	assign w_sub06_U_datain = ( (|r_sys_processing_methodID) ? r_sub06_U_datain : 32'h0 ) ;
	assign w_sub06_U_r_w = ( (|r_sys_processing_methodID) ? r_sub06_U_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 15'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_T_addr = ( (|r_sys_processing_methodID) ? r_sub15_T_addr : 15'sh0 ) ;
	assign w_sub15_T_datain = ( (|r_sys_processing_methodID) ? r_sub15_T_datain : 32'h0 ) ;
	assign w_sub15_T_r_w = ( (|r_sys_processing_methodID) ? r_sub15_T_r_w : 1'h0 ) ;
	assign w_sub15_V_addr = ( (|r_sys_processing_methodID) ? r_sub15_V_addr : 15'sh0 ) ;
	assign w_sub15_V_datain = ( (|r_sys_processing_methodID) ? r_sub15_V_datain : 32'h0 ) ;
	assign w_sub15_V_r_w = ( (|r_sys_processing_methodID) ? r_sub15_V_r_w : 1'h0 ) ;
	assign w_sub15_U_addr = ( (|r_sys_processing_methodID) ? r_sub15_U_addr : 15'sh0 ) ;
	assign w_sub15_U_datain = ( (|r_sys_processing_methodID) ? r_sub15_U_datain : 32'h0 ) ;
	assign w_sub15_U_r_w = ( (|r_sys_processing_methodID) ? r_sub15_U_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 15'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_T_addr = ( (|r_sys_processing_methodID) ? r_sub05_T_addr : 15'sh0 ) ;
	assign w_sub05_T_datain = ( (|r_sys_processing_methodID) ? r_sub05_T_datain : 32'h0 ) ;
	assign w_sub05_T_r_w = ( (|r_sys_processing_methodID) ? r_sub05_T_r_w : 1'h0 ) ;
	assign w_sub05_V_addr = ( (|r_sys_processing_methodID) ? r_sub05_V_addr : 15'sh0 ) ;
	assign w_sub05_V_datain = ( (|r_sys_processing_methodID) ? r_sub05_V_datain : 32'h0 ) ;
	assign w_sub05_V_r_w = ( (|r_sys_processing_methodID) ? r_sub05_V_r_w : 1'h0 ) ;
	assign w_sub05_U_addr = ( (|r_sys_processing_methodID) ? r_sub05_U_addr : 15'sh0 ) ;
	assign w_sub05_U_datain = ( (|r_sys_processing_methodID) ? r_sub05_U_datain : 32'h0 ) ;
	assign w_sub05_U_r_w = ( (|r_sys_processing_methodID) ? r_sub05_U_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 15'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_T_addr = ( (|r_sys_processing_methodID) ? r_sub04_T_addr : 15'sh0 ) ;
	assign w_sub04_T_datain = ( (|r_sys_processing_methodID) ? r_sub04_T_datain : 32'h0 ) ;
	assign w_sub04_T_r_w = ( (|r_sys_processing_methodID) ? r_sub04_T_r_w : 1'h0 ) ;
	assign w_sub04_V_addr = ( (|r_sys_processing_methodID) ? r_sub04_V_addr : 15'sh0 ) ;
	assign w_sub04_V_datain = ( (|r_sys_processing_methodID) ? r_sub04_V_datain : 32'h0 ) ;
	assign w_sub04_V_r_w = ( (|r_sys_processing_methodID) ? r_sub04_V_r_w : 1'h0 ) ;
	assign w_sub04_U_addr = ( (|r_sys_processing_methodID) ? r_sub04_U_addr : 15'sh0 ) ;
	assign w_sub04_U_datain = ( (|r_sys_processing_methodID) ? r_sub04_U_datain : 32'h0 ) ;
	assign w_sub04_U_r_w = ( (|r_sys_processing_methodID) ? r_sub04_U_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 15'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_T_addr = ( (|r_sys_processing_methodID) ? r_sub10_T_addr : 15'sh0 ) ;
	assign w_sub10_T_datain = ( (|r_sys_processing_methodID) ? r_sub10_T_datain : 32'h0 ) ;
	assign w_sub10_T_r_w = ( (|r_sys_processing_methodID) ? r_sub10_T_r_w : 1'h0 ) ;
	assign w_sub10_V_addr = ( (|r_sys_processing_methodID) ? r_sub10_V_addr : 15'sh0 ) ;
	assign w_sub10_V_datain = ( (|r_sys_processing_methodID) ? r_sub10_V_datain : 32'h0 ) ;
	assign w_sub10_V_r_w = ( (|r_sys_processing_methodID) ? r_sub10_V_r_w : 1'h0 ) ;
	assign w_sub10_U_addr = ( (|r_sys_processing_methodID) ? r_sub10_U_addr : 15'sh0 ) ;
	assign w_sub10_U_datain = ( (|r_sys_processing_methodID) ? r_sub10_U_datain : 32'h0 ) ;
	assign w_sub10_U_r_w = ( (|r_sys_processing_methodID) ? r_sub10_U_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 15'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000080;
	assign w_sys_tmp3 = 32'sh00000081;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'h3d000000;
	assign w_sys_tmp7 = 32'h3c000000;
	assign w_sys_tmp8 = 32'h3c03126f;
	assign w_sys_tmp9 = 32'h3d03126f;
	assign w_sys_tmp10 = 32'h3f03126f;
	assign w_sys_tmp11 = 32'h4103126f;
	assign w_sys_tmp12 = ( !w_sys_tmp13 );
	assign w_sys_tmp13 = (r_run_my_24 < r_run_k_20);
	assign w_sys_tmp14 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp15 = ( !w_sys_tmp16 );
	assign w_sys_tmp16 = (r_run_mx_23 < r_run_j_21);
	assign w_sys_tmp18 = w_ip_MultFloat_product_0;
	assign w_sys_tmp19 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp20 = (r_run_k_20 - w_sys_intOne);
	assign w_sys_tmp22 = (w_sys_tmp23 + r_run_k_20);
	assign w_sys_tmp23 = (r_run_j_21 * w_sys_tmp24);
	assign w_sys_tmp24 = 32'sh00000081;
	assign w_sys_tmp25 = 32'h0;
	assign w_sys_tmp27 = (w_sys_tmp28 + r_run_k_20);
	assign w_sys_tmp28 = (r_run_copy2_j_38 * w_sys_tmp24);
	assign w_sys_tmp32 = (w_sys_tmp33 + r_run_k_20);
	assign w_sys_tmp33 = (r_run_copy1_j_37 * w_sys_tmp24);
	assign w_sys_tmp36 = 32'h42200000;
	assign w_sys_tmp37 = w_sys_tmp18;
	assign w_sys_tmp38 = 32'h3f800000;
	assign w_sys_tmp41 = (w_sys_tmp42 + r_run_k_20);
	assign w_sys_tmp42 = (r_run_copy0_j_36 * w_sys_tmp24);
	assign w_sys_tmp45 = (r_run_copy0_j_36 + w_sys_intOne);
	assign w_sys_tmp46 = (r_run_copy1_j_37 + w_sys_intOne);
	assign w_sys_tmp47 = (r_run_copy2_j_38 + w_sys_intOne);
	assign w_sys_tmp48 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp128 = r_sys_tmp4_float;
	assign w_sys_tmp226 = ( !w_sys_tmp227 );
	assign w_sys_tmp227 = (w_sys_tmp228 < r_run_k_20);
	assign w_sys_tmp228 = 32'sh00000021;
	assign w_sys_tmp229 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp230 = ( !w_sys_tmp231 );
	assign w_sys_tmp231 = (w_sys_tmp232 < r_run_j_21);
	assign w_sys_tmp232 = 32'sh00000021;
	assign w_sys_tmp235 = (w_sys_tmp236 + r_run_k_20);
	assign w_sys_tmp236 = (r_run_j_21 * w_sys_tmp237);
	assign w_sys_tmp237 = 32'sh00000081;
	assign w_sys_tmp238 = w_fld_U_2_dataout_1;
	assign w_sys_tmp239 = (w_sys_tmp240 + r_run_k_20);
	assign w_sys_tmp240 = (r_run_copy4_j_43 * w_sys_tmp237);
	assign w_sys_tmp243 = (w_sys_tmp244 + r_run_k_20);
	assign w_sys_tmp244 = (r_run_copy3_j_42 * w_sys_tmp237);
	assign w_sys_tmp246 = w_fld_V_3_dataout_1;
	assign w_sys_tmp247 = (w_sys_tmp248 + r_run_k_20);
	assign w_sys_tmp248 = (r_run_copy2_j_41 * w_sys_tmp237);
	assign w_sys_tmp251 = (w_sys_tmp252 + r_run_k_20);
	assign w_sys_tmp252 = (r_run_copy1_j_40 * w_sys_tmp237);
	assign w_sys_tmp254 = w_fld_T_0_dataout_1;
	assign w_sys_tmp255 = (w_sys_tmp256 + r_run_k_20);
	assign w_sys_tmp256 = (r_run_copy0_j_39 * w_sys_tmp237);
	assign w_sys_tmp258 = (r_run_copy0_j_39 + w_sys_intOne);
	assign w_sys_tmp259 = (r_run_copy1_j_40 + w_sys_intOne);
	assign w_sys_tmp260 = (r_run_copy2_j_41 + w_sys_intOne);
	assign w_sys_tmp261 = (r_run_copy3_j_42 + w_sys_intOne);
	assign w_sys_tmp262 = (r_run_copy4_j_43 + w_sys_intOne);
	assign w_sys_tmp263 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp444 = 32'sh00000020;
	assign w_sys_tmp445 = ( !w_sys_tmp446 );
	assign w_sys_tmp446 = (w_sys_tmp447 < r_run_j_21);
	assign w_sys_tmp447 = 32'sh00000041;
	assign w_sys_tmp450 = (w_sys_tmp451 + r_run_k_20);
	assign w_sys_tmp451 = (r_run_j_21 * w_sys_tmp452);
	assign w_sys_tmp452 = 32'sh00000081;
	assign w_sys_tmp453 = w_fld_U_2_dataout_1;
	assign w_sys_tmp454 = (w_sys_tmp455 + r_run_k_20);
	assign w_sys_tmp455 = (r_run_copy4_j_48 * w_sys_tmp452);
	assign w_sys_tmp458 = (w_sys_tmp459 + r_run_k_20);
	assign w_sys_tmp459 = (r_run_copy3_j_47 * w_sys_tmp452);
	assign w_sys_tmp461 = w_fld_V_3_dataout_1;
	assign w_sys_tmp462 = (w_sys_tmp463 + r_run_k_20);
	assign w_sys_tmp463 = (r_run_copy2_j_46 * w_sys_tmp452);
	assign w_sys_tmp466 = (w_sys_tmp467 + r_run_k_20);
	assign w_sys_tmp467 = (r_run_copy1_j_45 * w_sys_tmp452);
	assign w_sys_tmp469 = w_fld_T_0_dataout_1;
	assign w_sys_tmp470 = (w_sys_tmp471 + r_run_k_20);
	assign w_sys_tmp471 = (r_run_copy0_j_44 * w_sys_tmp452);
	assign w_sys_tmp473 = (r_run_copy0_j_44 + w_sys_intOne);
	assign w_sys_tmp474 = (r_run_copy1_j_45 + w_sys_intOne);
	assign w_sys_tmp475 = (r_run_copy2_j_46 + w_sys_intOne);
	assign w_sys_tmp476 = (r_run_copy3_j_47 + w_sys_intOne);
	assign w_sys_tmp477 = (r_run_copy4_j_48 + w_sys_intOne);
	assign w_sys_tmp478 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp659 = 32'sh00000040;
	assign w_sys_tmp660 = ( !w_sys_tmp661 );
	assign w_sys_tmp661 = (w_sys_tmp662 < r_run_j_21);
	assign w_sys_tmp662 = 32'sh00000061;
	assign w_sys_tmp665 = (w_sys_tmp666 + r_run_k_20);
	assign w_sys_tmp666 = (r_run_j_21 * w_sys_tmp667);
	assign w_sys_tmp667 = 32'sh00000081;
	assign w_sys_tmp668 = w_fld_U_2_dataout_1;
	assign w_sys_tmp669 = (w_sys_tmp670 + r_run_k_20);
	assign w_sys_tmp670 = (r_run_copy4_j_53 * w_sys_tmp667);
	assign w_sys_tmp673 = (w_sys_tmp674 + r_run_k_20);
	assign w_sys_tmp674 = (r_run_copy3_j_52 * w_sys_tmp667);
	assign w_sys_tmp676 = w_fld_V_3_dataout_1;
	assign w_sys_tmp677 = (w_sys_tmp678 + r_run_k_20);
	assign w_sys_tmp678 = (r_run_copy2_j_51 * w_sys_tmp667);
	assign w_sys_tmp681 = (w_sys_tmp682 + r_run_k_20);
	assign w_sys_tmp682 = (r_run_copy1_j_50 * w_sys_tmp667);
	assign w_sys_tmp684 = w_fld_T_0_dataout_1;
	assign w_sys_tmp685 = (w_sys_tmp686 + r_run_k_20);
	assign w_sys_tmp686 = (r_run_copy0_j_49 * w_sys_tmp667);
	assign w_sys_tmp688 = (r_run_copy0_j_49 + w_sys_intOne);
	assign w_sys_tmp689 = (r_run_copy1_j_50 + w_sys_intOne);
	assign w_sys_tmp690 = (r_run_copy2_j_51 + w_sys_intOne);
	assign w_sys_tmp691 = (r_run_copy3_j_52 + w_sys_intOne);
	assign w_sys_tmp692 = (r_run_copy4_j_53 + w_sys_intOne);
	assign w_sys_tmp693 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp874 = 32'sh00000060;
	assign w_sys_tmp875 = ( !w_sys_tmp876 );
	assign w_sys_tmp876 = (w_sys_tmp877 < r_run_j_21);
	assign w_sys_tmp877 = 32'sh00000081;
	assign w_sys_tmp880 = (w_sys_tmp881 + r_run_k_20);
	assign w_sys_tmp881 = (r_run_j_21 * w_sys_tmp882);
	assign w_sys_tmp882 = 32'sh00000081;
	assign w_sys_tmp883 = w_fld_U_2_dataout_1;
	assign w_sys_tmp884 = (w_sys_tmp885 + r_run_k_20);
	assign w_sys_tmp885 = (r_run_copy4_j_58 * w_sys_tmp882);
	assign w_sys_tmp888 = (w_sys_tmp889 + r_run_k_20);
	assign w_sys_tmp889 = (r_run_copy3_j_57 * w_sys_tmp882);
	assign w_sys_tmp891 = w_fld_V_3_dataout_1;
	assign w_sys_tmp892 = (w_sys_tmp893 + r_run_k_20);
	assign w_sys_tmp893 = (r_run_copy2_j_56 * w_sys_tmp882);
	assign w_sys_tmp896 = (w_sys_tmp897 + r_run_k_20);
	assign w_sys_tmp897 = (r_run_copy1_j_55 * w_sys_tmp882);
	assign w_sys_tmp899 = w_fld_T_0_dataout_1;
	assign w_sys_tmp900 = (w_sys_tmp901 + r_run_k_20);
	assign w_sys_tmp901 = (r_run_copy0_j_54 * w_sys_tmp882);
	assign w_sys_tmp903 = (r_run_copy0_j_54 + w_sys_intOne);
	assign w_sys_tmp904 = (r_run_copy1_j_55 + w_sys_intOne);
	assign w_sys_tmp905 = (r_run_copy2_j_56 + w_sys_intOne);
	assign w_sys_tmp906 = (r_run_copy3_j_57 + w_sys_intOne);
	assign w_sys_tmp907 = (r_run_copy4_j_58 + w_sys_intOne);
	assign w_sys_tmp908 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp1089 = 32'sh00000020;
	assign w_sys_tmp1090 = ( !w_sys_tmp1091 );
	assign w_sys_tmp1091 = (w_sys_tmp1092 < r_run_k_20);
	assign w_sys_tmp1092 = 32'sh00000041;
	assign w_sys_tmp1093 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp1094 = ( !w_sys_tmp1095 );
	assign w_sys_tmp1095 = (w_sys_tmp1096 < r_run_j_21);
	assign w_sys_tmp1096 = 32'sh00000021;
	assign w_sys_tmp1099 = (w_sys_tmp1100 + r_run_k_20);
	assign w_sys_tmp1100 = (r_run_j_21 * w_sys_tmp1101);
	assign w_sys_tmp1101 = 32'sh00000081;
	assign w_sys_tmp1102 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1103 = (w_sys_tmp1104 + r_run_k_20);
	assign w_sys_tmp1104 = (r_run_copy4_j_63 * w_sys_tmp1101);
	assign w_sys_tmp1107 = (w_sys_tmp1108 + r_run_k_20);
	assign w_sys_tmp1108 = (r_run_copy3_j_62 * w_sys_tmp1101);
	assign w_sys_tmp1110 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1111 = (w_sys_tmp1112 + r_run_k_20);
	assign w_sys_tmp1112 = (r_run_copy2_j_61 * w_sys_tmp1101);
	assign w_sys_tmp1115 = (w_sys_tmp1116 + r_run_k_20);
	assign w_sys_tmp1116 = (r_run_copy1_j_60 * w_sys_tmp1101);
	assign w_sys_tmp1118 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1119 = (w_sys_tmp1120 + r_run_k_20);
	assign w_sys_tmp1120 = (r_run_copy0_j_59 * w_sys_tmp1101);
	assign w_sys_tmp1122 = (r_run_copy0_j_59 + w_sys_intOne);
	assign w_sys_tmp1123 = (r_run_copy1_j_60 + w_sys_intOne);
	assign w_sys_tmp1124 = (r_run_copy2_j_61 + w_sys_intOne);
	assign w_sys_tmp1125 = (r_run_copy3_j_62 + w_sys_intOne);
	assign w_sys_tmp1126 = (r_run_copy4_j_63 + w_sys_intOne);
	assign w_sys_tmp1127 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp1308 = 32'sh00000020;
	assign w_sys_tmp1309 = ( !w_sys_tmp1310 );
	assign w_sys_tmp1310 = (w_sys_tmp1311 < r_run_j_21);
	assign w_sys_tmp1311 = 32'sh00000041;
	assign w_sys_tmp1314 = (w_sys_tmp1315 + r_run_k_20);
	assign w_sys_tmp1315 = (r_run_j_21 * w_sys_tmp1316);
	assign w_sys_tmp1316 = 32'sh00000081;
	assign w_sys_tmp1317 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1318 = (w_sys_tmp1319 + r_run_k_20);
	assign w_sys_tmp1319 = (r_run_copy4_j_68 * w_sys_tmp1316);
	assign w_sys_tmp1322 = (w_sys_tmp1323 + r_run_k_20);
	assign w_sys_tmp1323 = (r_run_copy3_j_67 * w_sys_tmp1316);
	assign w_sys_tmp1325 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1326 = (w_sys_tmp1327 + r_run_k_20);
	assign w_sys_tmp1327 = (r_run_copy2_j_66 * w_sys_tmp1316);
	assign w_sys_tmp1330 = (w_sys_tmp1331 + r_run_k_20);
	assign w_sys_tmp1331 = (r_run_copy1_j_65 * w_sys_tmp1316);
	assign w_sys_tmp1333 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1334 = (w_sys_tmp1335 + r_run_k_20);
	assign w_sys_tmp1335 = (r_run_copy0_j_64 * w_sys_tmp1316);
	assign w_sys_tmp1337 = (r_run_copy0_j_64 + w_sys_intOne);
	assign w_sys_tmp1338 = (r_run_copy1_j_65 + w_sys_intOne);
	assign w_sys_tmp1339 = (r_run_copy2_j_66 + w_sys_intOne);
	assign w_sys_tmp1340 = (r_run_copy3_j_67 + w_sys_intOne);
	assign w_sys_tmp1341 = (r_run_copy4_j_68 + w_sys_intOne);
	assign w_sys_tmp1342 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp1523 = 32'sh00000040;
	assign w_sys_tmp1524 = ( !w_sys_tmp1525 );
	assign w_sys_tmp1525 = (w_sys_tmp1526 < r_run_j_21);
	assign w_sys_tmp1526 = 32'sh00000061;
	assign w_sys_tmp1529 = (w_sys_tmp1530 + r_run_k_20);
	assign w_sys_tmp1530 = (r_run_j_21 * w_sys_tmp1531);
	assign w_sys_tmp1531 = 32'sh00000081;
	assign w_sys_tmp1532 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1533 = (w_sys_tmp1534 + r_run_k_20);
	assign w_sys_tmp1534 = (r_run_copy4_j_73 * w_sys_tmp1531);
	assign w_sys_tmp1537 = (w_sys_tmp1538 + r_run_k_20);
	assign w_sys_tmp1538 = (r_run_copy3_j_72 * w_sys_tmp1531);
	assign w_sys_tmp1540 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1541 = (w_sys_tmp1542 + r_run_k_20);
	assign w_sys_tmp1542 = (r_run_copy2_j_71 * w_sys_tmp1531);
	assign w_sys_tmp1545 = (w_sys_tmp1546 + r_run_k_20);
	assign w_sys_tmp1546 = (r_run_copy1_j_70 * w_sys_tmp1531);
	assign w_sys_tmp1548 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1549 = (w_sys_tmp1550 + r_run_k_20);
	assign w_sys_tmp1550 = (r_run_copy0_j_69 * w_sys_tmp1531);
	assign w_sys_tmp1552 = (r_run_copy0_j_69 + w_sys_intOne);
	assign w_sys_tmp1553 = (r_run_copy1_j_70 + w_sys_intOne);
	assign w_sys_tmp1554 = (r_run_copy2_j_71 + w_sys_intOne);
	assign w_sys_tmp1555 = (r_run_copy3_j_72 + w_sys_intOne);
	assign w_sys_tmp1556 = (r_run_copy4_j_73 + w_sys_intOne);
	assign w_sys_tmp1557 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp1738 = 32'sh00000060;
	assign w_sys_tmp1739 = ( !w_sys_tmp1740 );
	assign w_sys_tmp1740 = (w_sys_tmp1741 < r_run_j_21);
	assign w_sys_tmp1741 = 32'sh00000081;
	assign w_sys_tmp1744 = (w_sys_tmp1745 + r_run_k_20);
	assign w_sys_tmp1745 = (r_run_j_21 * w_sys_tmp1746);
	assign w_sys_tmp1746 = 32'sh00000081;
	assign w_sys_tmp1747 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1748 = (w_sys_tmp1749 + r_run_k_20);
	assign w_sys_tmp1749 = (r_run_copy4_j_78 * w_sys_tmp1746);
	assign w_sys_tmp1752 = (w_sys_tmp1753 + r_run_k_20);
	assign w_sys_tmp1753 = (r_run_copy3_j_77 * w_sys_tmp1746);
	assign w_sys_tmp1755 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1756 = (w_sys_tmp1757 + r_run_k_20);
	assign w_sys_tmp1757 = (r_run_copy2_j_76 * w_sys_tmp1746);
	assign w_sys_tmp1760 = (w_sys_tmp1761 + r_run_k_20);
	assign w_sys_tmp1761 = (r_run_copy1_j_75 * w_sys_tmp1746);
	assign w_sys_tmp1763 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1764 = (w_sys_tmp1765 + r_run_k_20);
	assign w_sys_tmp1765 = (r_run_copy0_j_74 * w_sys_tmp1746);
	assign w_sys_tmp1767 = (r_run_copy0_j_74 + w_sys_intOne);
	assign w_sys_tmp1768 = (r_run_copy1_j_75 + w_sys_intOne);
	assign w_sys_tmp1769 = (r_run_copy2_j_76 + w_sys_intOne);
	assign w_sys_tmp1770 = (r_run_copy3_j_77 + w_sys_intOne);
	assign w_sys_tmp1771 = (r_run_copy4_j_78 + w_sys_intOne);
	assign w_sys_tmp1772 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp1953 = 32'sh00000040;
	assign w_sys_tmp1954 = ( !w_sys_tmp1955 );
	assign w_sys_tmp1955 = (w_sys_tmp1956 < r_run_k_20);
	assign w_sys_tmp1956 = 32'sh00000061;
	assign w_sys_tmp1957 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp1958 = ( !w_sys_tmp1959 );
	assign w_sys_tmp1959 = (w_sys_tmp1960 < r_run_j_21);
	assign w_sys_tmp1960 = 32'sh00000021;
	assign w_sys_tmp1963 = (w_sys_tmp1964 + r_run_k_20);
	assign w_sys_tmp1964 = (r_run_j_21 * w_sys_tmp1965);
	assign w_sys_tmp1965 = 32'sh00000081;
	assign w_sys_tmp1966 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1967 = (w_sys_tmp1968 + r_run_k_20);
	assign w_sys_tmp1968 = (r_run_copy4_j_83 * w_sys_tmp1965);
	assign w_sys_tmp1971 = (w_sys_tmp1972 + r_run_k_20);
	assign w_sys_tmp1972 = (r_run_copy3_j_82 * w_sys_tmp1965);
	assign w_sys_tmp1974 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1975 = (w_sys_tmp1976 + r_run_k_20);
	assign w_sys_tmp1976 = (r_run_copy2_j_81 * w_sys_tmp1965);
	assign w_sys_tmp1979 = (w_sys_tmp1980 + r_run_k_20);
	assign w_sys_tmp1980 = (r_run_copy1_j_80 * w_sys_tmp1965);
	assign w_sys_tmp1982 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1983 = (w_sys_tmp1984 + r_run_k_20);
	assign w_sys_tmp1984 = (r_run_copy0_j_79 * w_sys_tmp1965);
	assign w_sys_tmp1986 = (r_run_copy0_j_79 + w_sys_intOne);
	assign w_sys_tmp1987 = (r_run_copy1_j_80 + w_sys_intOne);
	assign w_sys_tmp1988 = (r_run_copy2_j_81 + w_sys_intOne);
	assign w_sys_tmp1989 = (r_run_copy3_j_82 + w_sys_intOne);
	assign w_sys_tmp1990 = (r_run_copy4_j_83 + w_sys_intOne);
	assign w_sys_tmp1991 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp2172 = 32'sh00000020;
	assign w_sys_tmp2173 = ( !w_sys_tmp2174 );
	assign w_sys_tmp2174 = (w_sys_tmp2175 < r_run_j_21);
	assign w_sys_tmp2175 = 32'sh00000041;
	assign w_sys_tmp2178 = (w_sys_tmp2179 + r_run_k_20);
	assign w_sys_tmp2179 = (r_run_j_21 * w_sys_tmp2180);
	assign w_sys_tmp2180 = 32'sh00000081;
	assign w_sys_tmp2181 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2182 = (w_sys_tmp2183 + r_run_k_20);
	assign w_sys_tmp2183 = (r_run_copy4_j_88 * w_sys_tmp2180);
	assign w_sys_tmp2186 = (w_sys_tmp2187 + r_run_k_20);
	assign w_sys_tmp2187 = (r_run_copy3_j_87 * w_sys_tmp2180);
	assign w_sys_tmp2189 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2190 = (w_sys_tmp2191 + r_run_k_20);
	assign w_sys_tmp2191 = (r_run_copy2_j_86 * w_sys_tmp2180);
	assign w_sys_tmp2194 = (w_sys_tmp2195 + r_run_k_20);
	assign w_sys_tmp2195 = (r_run_copy1_j_85 * w_sys_tmp2180);
	assign w_sys_tmp2197 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2198 = (w_sys_tmp2199 + r_run_k_20);
	assign w_sys_tmp2199 = (r_run_copy0_j_84 * w_sys_tmp2180);
	assign w_sys_tmp2201 = (r_run_copy0_j_84 + w_sys_intOne);
	assign w_sys_tmp2202 = (r_run_copy1_j_85 + w_sys_intOne);
	assign w_sys_tmp2203 = (r_run_copy2_j_86 + w_sys_intOne);
	assign w_sys_tmp2204 = (r_run_copy3_j_87 + w_sys_intOne);
	assign w_sys_tmp2205 = (r_run_copy4_j_88 + w_sys_intOne);
	assign w_sys_tmp2206 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp2387 = 32'sh00000040;
	assign w_sys_tmp2388 = ( !w_sys_tmp2389 );
	assign w_sys_tmp2389 = (w_sys_tmp2390 < r_run_j_21);
	assign w_sys_tmp2390 = 32'sh00000061;
	assign w_sys_tmp2393 = (w_sys_tmp2394 + r_run_k_20);
	assign w_sys_tmp2394 = (r_run_j_21 * w_sys_tmp2395);
	assign w_sys_tmp2395 = 32'sh00000081;
	assign w_sys_tmp2396 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2397 = (w_sys_tmp2398 + r_run_k_20);
	assign w_sys_tmp2398 = (r_run_copy4_j_93 * w_sys_tmp2395);
	assign w_sys_tmp2401 = (w_sys_tmp2402 + r_run_k_20);
	assign w_sys_tmp2402 = (r_run_copy3_j_92 * w_sys_tmp2395);
	assign w_sys_tmp2404 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2405 = (w_sys_tmp2406 + r_run_k_20);
	assign w_sys_tmp2406 = (r_run_copy2_j_91 * w_sys_tmp2395);
	assign w_sys_tmp2409 = (w_sys_tmp2410 + r_run_k_20);
	assign w_sys_tmp2410 = (r_run_copy1_j_90 * w_sys_tmp2395);
	assign w_sys_tmp2412 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2413 = (w_sys_tmp2414 + r_run_k_20);
	assign w_sys_tmp2414 = (r_run_copy0_j_89 * w_sys_tmp2395);
	assign w_sys_tmp2416 = (r_run_copy0_j_89 + w_sys_intOne);
	assign w_sys_tmp2417 = (r_run_copy1_j_90 + w_sys_intOne);
	assign w_sys_tmp2418 = (r_run_copy2_j_91 + w_sys_intOne);
	assign w_sys_tmp2419 = (r_run_copy3_j_92 + w_sys_intOne);
	assign w_sys_tmp2420 = (r_run_copy4_j_93 + w_sys_intOne);
	assign w_sys_tmp2421 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp2602 = 32'sh00000060;
	assign w_sys_tmp2603 = ( !w_sys_tmp2604 );
	assign w_sys_tmp2604 = (w_sys_tmp2605 < r_run_j_21);
	assign w_sys_tmp2605 = 32'sh00000081;
	assign w_sys_tmp2608 = (w_sys_tmp2609 + r_run_k_20);
	assign w_sys_tmp2609 = (r_run_j_21 * w_sys_tmp2610);
	assign w_sys_tmp2610 = 32'sh00000081;
	assign w_sys_tmp2611 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2612 = (w_sys_tmp2613 + r_run_k_20);
	assign w_sys_tmp2613 = (r_run_copy4_j_98 * w_sys_tmp2610);
	assign w_sys_tmp2616 = (w_sys_tmp2617 + r_run_k_20);
	assign w_sys_tmp2617 = (r_run_copy3_j_97 * w_sys_tmp2610);
	assign w_sys_tmp2619 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2620 = (w_sys_tmp2621 + r_run_k_20);
	assign w_sys_tmp2621 = (r_run_copy2_j_96 * w_sys_tmp2610);
	assign w_sys_tmp2624 = (w_sys_tmp2625 + r_run_k_20);
	assign w_sys_tmp2625 = (r_run_copy1_j_95 * w_sys_tmp2610);
	assign w_sys_tmp2627 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2628 = (w_sys_tmp2629 + r_run_k_20);
	assign w_sys_tmp2629 = (r_run_copy0_j_94 * w_sys_tmp2610);
	assign w_sys_tmp2631 = (r_run_copy0_j_94 + w_sys_intOne);
	assign w_sys_tmp2632 = (r_run_copy1_j_95 + w_sys_intOne);
	assign w_sys_tmp2633 = (r_run_copy2_j_96 + w_sys_intOne);
	assign w_sys_tmp2634 = (r_run_copy3_j_97 + w_sys_intOne);
	assign w_sys_tmp2635 = (r_run_copy4_j_98 + w_sys_intOne);
	assign w_sys_tmp2636 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp2817 = 32'sh00000060;
	assign w_sys_tmp2818 = ( !w_sys_tmp2819 );
	assign w_sys_tmp2819 = (w_sys_tmp2820 < r_run_k_20);
	assign w_sys_tmp2820 = 32'sh00000081;
	assign w_sys_tmp2821 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp2822 = ( !w_sys_tmp2823 );
	assign w_sys_tmp2823 = (w_sys_tmp2824 < r_run_j_21);
	assign w_sys_tmp2824 = 32'sh00000021;
	assign w_sys_tmp2827 = (w_sys_tmp2828 + r_run_k_20);
	assign w_sys_tmp2828 = (r_run_j_21 * w_sys_tmp2829);
	assign w_sys_tmp2829 = 32'sh00000081;
	assign w_sys_tmp2830 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2831 = (w_sys_tmp2832 + r_run_k_20);
	assign w_sys_tmp2832 = (r_run_copy4_j_103 * w_sys_tmp2829);
	assign w_sys_tmp2835 = (w_sys_tmp2836 + r_run_k_20);
	assign w_sys_tmp2836 = (r_run_copy3_j_102 * w_sys_tmp2829);
	assign w_sys_tmp2838 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2839 = (w_sys_tmp2840 + r_run_k_20);
	assign w_sys_tmp2840 = (r_run_copy2_j_101 * w_sys_tmp2829);
	assign w_sys_tmp2843 = (w_sys_tmp2844 + r_run_k_20);
	assign w_sys_tmp2844 = (r_run_copy1_j_100 * w_sys_tmp2829);
	assign w_sys_tmp2846 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2847 = (w_sys_tmp2848 + r_run_k_20);
	assign w_sys_tmp2848 = (r_run_copy0_j_99 * w_sys_tmp2829);
	assign w_sys_tmp2850 = (r_run_copy0_j_99 + w_sys_intOne);
	assign w_sys_tmp2851 = (r_run_copy1_j_100 + w_sys_intOne);
	assign w_sys_tmp2852 = (r_run_copy2_j_101 + w_sys_intOne);
	assign w_sys_tmp2853 = (r_run_copy3_j_102 + w_sys_intOne);
	assign w_sys_tmp2854 = (r_run_copy4_j_103 + w_sys_intOne);
	assign w_sys_tmp2855 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp3036 = 32'sh00000020;
	assign w_sys_tmp3037 = ( !w_sys_tmp3038 );
	assign w_sys_tmp3038 = (w_sys_tmp3039 < r_run_j_21);
	assign w_sys_tmp3039 = 32'sh00000041;
	assign w_sys_tmp3042 = (w_sys_tmp3043 + r_run_k_20);
	assign w_sys_tmp3043 = (r_run_j_21 * w_sys_tmp3044);
	assign w_sys_tmp3044 = 32'sh00000081;
	assign w_sys_tmp3045 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3046 = (w_sys_tmp3047 + r_run_k_20);
	assign w_sys_tmp3047 = (r_run_copy4_j_108 * w_sys_tmp3044);
	assign w_sys_tmp3050 = (w_sys_tmp3051 + r_run_k_20);
	assign w_sys_tmp3051 = (r_run_copy3_j_107 * w_sys_tmp3044);
	assign w_sys_tmp3053 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3054 = (w_sys_tmp3055 + r_run_k_20);
	assign w_sys_tmp3055 = (r_run_copy2_j_106 * w_sys_tmp3044);
	assign w_sys_tmp3058 = (w_sys_tmp3059 + r_run_k_20);
	assign w_sys_tmp3059 = (r_run_copy1_j_105 * w_sys_tmp3044);
	assign w_sys_tmp3061 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3062 = (w_sys_tmp3063 + r_run_k_20);
	assign w_sys_tmp3063 = (r_run_copy0_j_104 * w_sys_tmp3044);
	assign w_sys_tmp3065 = (r_run_copy0_j_104 + w_sys_intOne);
	assign w_sys_tmp3066 = (r_run_copy1_j_105 + w_sys_intOne);
	assign w_sys_tmp3067 = (r_run_copy2_j_106 + w_sys_intOne);
	assign w_sys_tmp3068 = (r_run_copy3_j_107 + w_sys_intOne);
	assign w_sys_tmp3069 = (r_run_copy4_j_108 + w_sys_intOne);
	assign w_sys_tmp3070 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp3251 = 32'sh00000040;
	assign w_sys_tmp3252 = ( !w_sys_tmp3253 );
	assign w_sys_tmp3253 = (w_sys_tmp3254 < r_run_j_21);
	assign w_sys_tmp3254 = 32'sh00000061;
	assign w_sys_tmp3257 = (w_sys_tmp3258 + r_run_k_20);
	assign w_sys_tmp3258 = (r_run_j_21 * w_sys_tmp3259);
	assign w_sys_tmp3259 = 32'sh00000081;
	assign w_sys_tmp3260 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3261 = (w_sys_tmp3262 + r_run_k_20);
	assign w_sys_tmp3262 = (r_run_copy4_j_113 * w_sys_tmp3259);
	assign w_sys_tmp3265 = (w_sys_tmp3266 + r_run_k_20);
	assign w_sys_tmp3266 = (r_run_copy3_j_112 * w_sys_tmp3259);
	assign w_sys_tmp3268 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3269 = (w_sys_tmp3270 + r_run_k_20);
	assign w_sys_tmp3270 = (r_run_copy2_j_111 * w_sys_tmp3259);
	assign w_sys_tmp3273 = (w_sys_tmp3274 + r_run_k_20);
	assign w_sys_tmp3274 = (r_run_copy1_j_110 * w_sys_tmp3259);
	assign w_sys_tmp3276 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3277 = (w_sys_tmp3278 + r_run_k_20);
	assign w_sys_tmp3278 = (r_run_copy0_j_109 * w_sys_tmp3259);
	assign w_sys_tmp3280 = (r_run_copy0_j_109 + w_sys_intOne);
	assign w_sys_tmp3281 = (r_run_copy1_j_110 + w_sys_intOne);
	assign w_sys_tmp3282 = (r_run_copy2_j_111 + w_sys_intOne);
	assign w_sys_tmp3283 = (r_run_copy3_j_112 + w_sys_intOne);
	assign w_sys_tmp3284 = (r_run_copy4_j_113 + w_sys_intOne);
	assign w_sys_tmp3285 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp3466 = 32'sh00000060;
	assign w_sys_tmp3467 = ( !w_sys_tmp3468 );
	assign w_sys_tmp3468 = (w_sys_tmp3469 < r_run_j_21);
	assign w_sys_tmp3469 = 32'sh00000081;
	assign w_sys_tmp3472 = (w_sys_tmp3473 + r_run_k_20);
	assign w_sys_tmp3473 = (r_run_j_21 * w_sys_tmp3474);
	assign w_sys_tmp3474 = 32'sh00000081;
	assign w_sys_tmp3475 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3476 = (w_sys_tmp3477 + r_run_k_20);
	assign w_sys_tmp3477 = (r_run_copy4_j_118 * w_sys_tmp3474);
	assign w_sys_tmp3480 = (w_sys_tmp3481 + r_run_k_20);
	assign w_sys_tmp3481 = (r_run_copy3_j_117 * w_sys_tmp3474);
	assign w_sys_tmp3483 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3484 = (w_sys_tmp3485 + r_run_k_20);
	assign w_sys_tmp3485 = (r_run_copy2_j_116 * w_sys_tmp3474);
	assign w_sys_tmp3488 = (w_sys_tmp3489 + r_run_k_20);
	assign w_sys_tmp3489 = (r_run_copy1_j_115 * w_sys_tmp3474);
	assign w_sys_tmp3491 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3492 = (w_sys_tmp3493 + r_run_k_20);
	assign w_sys_tmp3493 = (r_run_copy0_j_114 * w_sys_tmp3474);
	assign w_sys_tmp3495 = (r_run_copy0_j_114 + w_sys_intOne);
	assign w_sys_tmp3496 = (r_run_copy1_j_115 + w_sys_intOne);
	assign w_sys_tmp3497 = (r_run_copy2_j_116 + w_sys_intOne);
	assign w_sys_tmp3498 = (r_run_copy3_j_117 + w_sys_intOne);
	assign w_sys_tmp3499 = (r_run_copy4_j_118 + w_sys_intOne);
	assign w_sys_tmp3500 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp3681 = ( !w_sys_tmp3682 );
	assign w_sys_tmp3682 = (r_run_nlast_35 < r_run_n_22);
	assign w_sys_tmp3683 = (r_run_n_22 + w_sys_intOne);
	assign w_sys_tmp3684 = 32'sh00000002;
	assign w_sys_tmp3685 = ( !w_sys_tmp3686 );
	assign w_sys_tmp3686 = (w_sys_tmp3687 < r_run_k_20);
	assign w_sys_tmp3687 = 32'sh00000020;
	assign w_sys_tmp3690 = (w_sys_tmp3691 + r_run_k_20);
	assign w_sys_tmp3691 = 32'sh000010a1;
	assign w_sys_tmp3692 = w_sub04_result_dataout;
	assign w_sys_tmp3696 = (w_sys_tmp3697 + r_run_k_20);
	assign w_sys_tmp3697 = 32'sh00001020;
	assign w_sys_tmp3698 = w_sub00_result_dataout;
	assign w_sys_tmp3702 = (w_sys_tmp3703 + r_run_k_20);
	assign w_sys_tmp3703 = 32'sh000020c1;
	assign w_sys_tmp3707 = (w_sys_tmp3708 + r_run_k_20);
	assign w_sys_tmp3708 = 32'sh00002040;
	assign w_sys_tmp3713 = (w_sys_tmp3714 + r_run_k_20);
	assign w_sys_tmp3714 = 32'sh000030e1;
	assign w_sys_tmp3718 = (w_sys_tmp3719 + r_run_k_20);
	assign w_sys_tmp3719 = 32'sh00003060;
	assign w_sys_tmp3720 = w_sub08_result_dataout;
	assign w_sys_tmp3723 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp3724 = 32'sh00000021;
	assign w_sys_tmp3725 = ( !w_sys_tmp3726 );
	assign w_sys_tmp3726 = (w_sys_tmp3727 < r_run_k_20);
	assign w_sys_tmp3727 = 32'sh00000040;
	assign w_sys_tmp3730 = (w_sys_tmp3731 + r_run_k_20);
	assign w_sys_tmp3731 = 32'sh000010a1;
	assign w_sys_tmp3732 = w_sub05_result_dataout;
	assign w_sys_tmp3736 = (w_sys_tmp3737 + r_run_k_20);
	assign w_sys_tmp3737 = 32'sh00001020;
	assign w_sys_tmp3738 = w_sub01_result_dataout;
	assign w_sys_tmp3742 = (w_sys_tmp3743 + r_run_k_20);
	assign w_sys_tmp3743 = 32'sh000020c1;
	assign w_sys_tmp3747 = (w_sys_tmp3748 + r_run_k_20);
	assign w_sys_tmp3748 = 32'sh00002040;
	assign w_sys_tmp3753 = (w_sys_tmp3754 + r_run_k_20);
	assign w_sys_tmp3754 = 32'sh000030e1;
	assign w_sys_tmp3758 = (w_sys_tmp3759 + r_run_k_20);
	assign w_sys_tmp3759 = 32'sh00003060;
	assign w_sys_tmp3760 = w_sub09_result_dataout;
	assign w_sys_tmp3763 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp3764 = 32'sh00000041;
	assign w_sys_tmp3765 = ( !w_sys_tmp3766 );
	assign w_sys_tmp3766 = (w_sys_tmp3767 < r_run_k_20);
	assign w_sys_tmp3767 = 32'sh00000060;
	assign w_sys_tmp3770 = (w_sys_tmp3771 + r_run_k_20);
	assign w_sys_tmp3771 = 32'sh000010a1;
	assign w_sys_tmp3772 = w_sub06_result_dataout;
	assign w_sys_tmp3776 = (w_sys_tmp3777 + r_run_k_20);
	assign w_sys_tmp3777 = 32'sh00001020;
	assign w_sys_tmp3778 = w_sub02_result_dataout;
	assign w_sys_tmp3782 = (w_sys_tmp3783 + r_run_k_20);
	assign w_sys_tmp3783 = 32'sh000020c1;
	assign w_sys_tmp3787 = (w_sys_tmp3788 + r_run_k_20);
	assign w_sys_tmp3788 = 32'sh00002040;
	assign w_sys_tmp3793 = (w_sys_tmp3794 + r_run_k_20);
	assign w_sys_tmp3794 = 32'sh000030e1;
	assign w_sys_tmp3798 = (w_sys_tmp3799 + r_run_k_20);
	assign w_sys_tmp3799 = 32'sh00003060;
	assign w_sys_tmp3800 = w_sub10_result_dataout;
	assign w_sys_tmp3803 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp3804 = 32'sh00000061;
	assign w_sys_tmp3805 = ( !w_sys_tmp3806 );
	assign w_sys_tmp3806 = (w_sys_tmp3807 < r_run_k_20);
	assign w_sys_tmp3807 = 32'sh00000080;
	assign w_sys_tmp3810 = (w_sys_tmp3811 + r_run_k_20);
	assign w_sys_tmp3811 = 32'sh000010a1;
	assign w_sys_tmp3812 = w_sub07_result_dataout;
	assign w_sys_tmp3816 = (w_sys_tmp3817 + r_run_k_20);
	assign w_sys_tmp3817 = 32'sh00001020;
	assign w_sys_tmp3818 = w_sub03_result_dataout;
	assign w_sys_tmp3822 = (w_sys_tmp3823 + r_run_k_20);
	assign w_sys_tmp3823 = 32'sh000020c1;
	assign w_sys_tmp3827 = (w_sys_tmp3828 + r_run_k_20);
	assign w_sys_tmp3828 = 32'sh00002040;
	assign w_sys_tmp3833 = (w_sys_tmp3834 + r_run_k_20);
	assign w_sys_tmp3834 = 32'sh000030e1;
	assign w_sys_tmp3838 = (w_sys_tmp3839 + r_run_k_20);
	assign w_sys_tmp3839 = 32'sh00003060;
	assign w_sys_tmp3840 = w_sub11_result_dataout;
	assign w_sys_tmp3843 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp3844 = 32'sh00000002;
	assign w_sys_tmp3845 = ( !w_sys_tmp3846 );
	assign w_sys_tmp3846 = (w_sys_tmp3847 < r_run_j_21);
	assign w_sys_tmp3847 = 32'sh00000020;
	assign w_sys_tmp3850 = (w_sys_tmp3851 + w_sys_tmp3853);
	assign w_sys_tmp3851 = (r_run_j_21 * w_sys_tmp3852);
	assign w_sys_tmp3852 = 32'sh00000081;
	assign w_sys_tmp3853 = 32'sh00000021;
	assign w_sys_tmp3854 = w_sub01_result_dataout;
	assign w_sys_tmp3855 = (w_sys_tmp3856 + w_sys_tmp3853);
	assign w_sys_tmp3856 = (r_run_copy10_j_129 * w_sys_tmp3852);
	assign w_sys_tmp3860 = (w_sys_tmp3861 + w_sys_tmp3863);
	assign w_sys_tmp3861 = (r_run_copy9_j_128 * w_sys_tmp3852);
	assign w_sys_tmp3863 = 32'sh00000020;
	assign w_sys_tmp3864 = w_sub00_result_dataout;
	assign w_sys_tmp3865 = (w_sys_tmp3866 + w_sys_tmp3863);
	assign w_sys_tmp3866 = (r_run_copy8_j_127 * w_sys_tmp3852);
	assign w_sys_tmp3870 = (w_sys_tmp3871 + w_sys_tmp3873);
	assign w_sys_tmp3871 = (r_run_copy7_j_126 * w_sys_tmp3852);
	assign w_sys_tmp3873 = 32'sh00000041;
	assign w_sys_tmp3874 = (w_sys_tmp3875 + w_sys_tmp3873);
	assign w_sys_tmp3875 = (r_run_copy6_j_125 * w_sys_tmp3852);
	assign w_sys_tmp3879 = (w_sys_tmp3880 + w_sys_tmp3882);
	assign w_sys_tmp3880 = (r_run_copy5_j_124 * w_sys_tmp3852);
	assign w_sys_tmp3882 = 32'sh00000040;
	assign w_sys_tmp3884 = (w_sys_tmp3885 + w_sys_tmp3882);
	assign w_sys_tmp3885 = (r_run_copy4_j_123 * w_sys_tmp3852);
	assign w_sys_tmp3889 = (w_sys_tmp3890 + w_sys_tmp3892);
	assign w_sys_tmp3890 = (r_run_copy3_j_122 * w_sys_tmp3852);
	assign w_sys_tmp3892 = 32'sh00000061;
	assign w_sys_tmp3893 = (w_sys_tmp3894 + w_sys_tmp3892);
	assign w_sys_tmp3894 = (r_run_copy2_j_121 * w_sys_tmp3852);
	assign w_sys_tmp3898 = (w_sys_tmp3899 + w_sys_tmp3901);
	assign w_sys_tmp3899 = (r_run_copy1_j_120 * w_sys_tmp3852);
	assign w_sys_tmp3901 = 32'sh00000060;
	assign w_sys_tmp3902 = w_sub02_result_dataout;
	assign w_sys_tmp3903 = (w_sys_tmp3904 + w_sys_tmp3901);
	assign w_sys_tmp3904 = (r_run_copy0_j_119 * w_sys_tmp3852);
	assign w_sys_tmp3907 = (r_run_copy0_j_119 + w_sys_intOne);
	assign w_sys_tmp3908 = (r_run_copy1_j_120 + w_sys_intOne);
	assign w_sys_tmp3909 = (r_run_copy2_j_121 + w_sys_intOne);
	assign w_sys_tmp3910 = (r_run_copy3_j_122 + w_sys_intOne);
	assign w_sys_tmp3911 = (r_run_copy4_j_123 + w_sys_intOne);
	assign w_sys_tmp3912 = (r_run_copy5_j_124 + w_sys_intOne);
	assign w_sys_tmp3913 = (r_run_copy6_j_125 + w_sys_intOne);
	assign w_sys_tmp3914 = (r_run_copy7_j_126 + w_sys_intOne);
	assign w_sys_tmp3915 = (r_run_copy8_j_127 + w_sys_intOne);
	assign w_sys_tmp3916 = (r_run_copy9_j_128 + w_sys_intOne);
	assign w_sys_tmp3917 = (r_run_copy10_j_129 + w_sys_intOne);
	assign w_sys_tmp3918 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp4345 = 32'sh00000021;
	assign w_sys_tmp4346 = ( !w_sys_tmp4347 );
	assign w_sys_tmp4347 = (w_sys_tmp4348 < r_run_j_21);
	assign w_sys_tmp4348 = 32'sh00000040;
	assign w_sys_tmp4351 = (w_sys_tmp4352 + w_sys_tmp4354);
	assign w_sys_tmp4352 = (r_run_j_21 * w_sys_tmp4353);
	assign w_sys_tmp4353 = 32'sh00000081;
	assign w_sys_tmp4354 = 32'sh00000021;
	assign w_sys_tmp4355 = w_sub05_result_dataout;
	assign w_sys_tmp4356 = (w_sys_tmp4357 + w_sys_tmp4354);
	assign w_sys_tmp4357 = (r_run_copy10_j_140 * w_sys_tmp4353);
	assign w_sys_tmp4361 = (w_sys_tmp4362 + w_sys_tmp4364);
	assign w_sys_tmp4362 = (r_run_copy9_j_139 * w_sys_tmp4353);
	assign w_sys_tmp4364 = 32'sh00000020;
	assign w_sys_tmp4365 = w_sub04_result_dataout;
	assign w_sys_tmp4366 = (w_sys_tmp4367 + w_sys_tmp4364);
	assign w_sys_tmp4367 = (r_run_copy8_j_138 * w_sys_tmp4353);
	assign w_sys_tmp4371 = (w_sys_tmp4372 + w_sys_tmp4374);
	assign w_sys_tmp4372 = (r_run_copy7_j_137 * w_sys_tmp4353);
	assign w_sys_tmp4374 = 32'sh00000041;
	assign w_sys_tmp4375 = (w_sys_tmp4376 + w_sys_tmp4374);
	assign w_sys_tmp4376 = (r_run_copy6_j_136 * w_sys_tmp4353);
	assign w_sys_tmp4380 = (w_sys_tmp4381 + w_sys_tmp4383);
	assign w_sys_tmp4381 = (r_run_copy5_j_135 * w_sys_tmp4353);
	assign w_sys_tmp4383 = 32'sh00000040;
	assign w_sys_tmp4385 = (w_sys_tmp4386 + w_sys_tmp4383);
	assign w_sys_tmp4386 = (r_run_copy4_j_134 * w_sys_tmp4353);
	assign w_sys_tmp4390 = (w_sys_tmp4391 + w_sys_tmp4393);
	assign w_sys_tmp4391 = (r_run_copy3_j_133 * w_sys_tmp4353);
	assign w_sys_tmp4393 = 32'sh00000061;
	assign w_sys_tmp4394 = (w_sys_tmp4395 + w_sys_tmp4393);
	assign w_sys_tmp4395 = (r_run_copy2_j_132 * w_sys_tmp4353);
	assign w_sys_tmp4399 = (w_sys_tmp4400 + w_sys_tmp4402);
	assign w_sys_tmp4400 = (r_run_copy1_j_131 * w_sys_tmp4353);
	assign w_sys_tmp4402 = 32'sh00000060;
	assign w_sys_tmp4403 = w_sub06_result_dataout;
	assign w_sys_tmp4404 = (w_sys_tmp4405 + w_sys_tmp4402);
	assign w_sys_tmp4405 = (r_run_copy0_j_130 * w_sys_tmp4353);
	assign w_sys_tmp4408 = (r_run_copy0_j_130 + w_sys_intOne);
	assign w_sys_tmp4409 = (r_run_copy1_j_131 + w_sys_intOne);
	assign w_sys_tmp4410 = (r_run_copy2_j_132 + w_sys_intOne);
	assign w_sys_tmp4411 = (r_run_copy3_j_133 + w_sys_intOne);
	assign w_sys_tmp4412 = (r_run_copy4_j_134 + w_sys_intOne);
	assign w_sys_tmp4413 = (r_run_copy5_j_135 + w_sys_intOne);
	assign w_sys_tmp4414 = (r_run_copy6_j_136 + w_sys_intOne);
	assign w_sys_tmp4415 = (r_run_copy7_j_137 + w_sys_intOne);
	assign w_sys_tmp4416 = (r_run_copy8_j_138 + w_sys_intOne);
	assign w_sys_tmp4417 = (r_run_copy9_j_139 + w_sys_intOne);
	assign w_sys_tmp4418 = (r_run_copy10_j_140 + w_sys_intOne);
	assign w_sys_tmp4419 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp4846 = 32'sh00000041;
	assign w_sys_tmp4847 = ( !w_sys_tmp4848 );
	assign w_sys_tmp4848 = (w_sys_tmp4849 < r_run_j_21);
	assign w_sys_tmp4849 = 32'sh00000060;
	assign w_sys_tmp4852 = (w_sys_tmp4853 + w_sys_tmp4855);
	assign w_sys_tmp4853 = (r_run_j_21 * w_sys_tmp4854);
	assign w_sys_tmp4854 = 32'sh00000081;
	assign w_sys_tmp4855 = 32'sh00000021;
	assign w_sys_tmp4856 = w_sub09_result_dataout;
	assign w_sys_tmp4857 = (w_sys_tmp4858 + w_sys_tmp4855);
	assign w_sys_tmp4858 = (r_run_copy10_j_151 * w_sys_tmp4854);
	assign w_sys_tmp4862 = (w_sys_tmp4863 + w_sys_tmp4865);
	assign w_sys_tmp4863 = (r_run_copy9_j_150 * w_sys_tmp4854);
	assign w_sys_tmp4865 = 32'sh00000020;
	assign w_sys_tmp4866 = w_sub08_result_dataout;
	assign w_sys_tmp4867 = (w_sys_tmp4868 + w_sys_tmp4865);
	assign w_sys_tmp4868 = (r_run_copy8_j_149 * w_sys_tmp4854);
	assign w_sys_tmp4872 = (w_sys_tmp4873 + w_sys_tmp4875);
	assign w_sys_tmp4873 = (r_run_copy7_j_148 * w_sys_tmp4854);
	assign w_sys_tmp4875 = 32'sh00000041;
	assign w_sys_tmp4876 = (w_sys_tmp4877 + w_sys_tmp4875);
	assign w_sys_tmp4877 = (r_run_copy6_j_147 * w_sys_tmp4854);
	assign w_sys_tmp4881 = (w_sys_tmp4882 + w_sys_tmp4884);
	assign w_sys_tmp4882 = (r_run_copy5_j_146 * w_sys_tmp4854);
	assign w_sys_tmp4884 = 32'sh00000040;
	assign w_sys_tmp4886 = (w_sys_tmp4887 + w_sys_tmp4884);
	assign w_sys_tmp4887 = (r_run_copy4_j_145 * w_sys_tmp4854);
	assign w_sys_tmp4891 = (w_sys_tmp4892 + w_sys_tmp4894);
	assign w_sys_tmp4892 = (r_run_copy3_j_144 * w_sys_tmp4854);
	assign w_sys_tmp4894 = 32'sh00000061;
	assign w_sys_tmp4895 = (w_sys_tmp4896 + w_sys_tmp4894);
	assign w_sys_tmp4896 = (r_run_copy2_j_143 * w_sys_tmp4854);
	assign w_sys_tmp4900 = (w_sys_tmp4901 + w_sys_tmp4903);
	assign w_sys_tmp4901 = (r_run_copy1_j_142 * w_sys_tmp4854);
	assign w_sys_tmp4903 = 32'sh00000060;
	assign w_sys_tmp4904 = w_sub10_result_dataout;
	assign w_sys_tmp4905 = (w_sys_tmp4906 + w_sys_tmp4903);
	assign w_sys_tmp4906 = (r_run_copy0_j_141 * w_sys_tmp4854);
	assign w_sys_tmp4909 = (r_run_copy0_j_141 + w_sys_intOne);
	assign w_sys_tmp4910 = (r_run_copy1_j_142 + w_sys_intOne);
	assign w_sys_tmp4911 = (r_run_copy2_j_143 + w_sys_intOne);
	assign w_sys_tmp4912 = (r_run_copy3_j_144 + w_sys_intOne);
	assign w_sys_tmp4913 = (r_run_copy4_j_145 + w_sys_intOne);
	assign w_sys_tmp4914 = (r_run_copy5_j_146 + w_sys_intOne);
	assign w_sys_tmp4915 = (r_run_copy6_j_147 + w_sys_intOne);
	assign w_sys_tmp4916 = (r_run_copy7_j_148 + w_sys_intOne);
	assign w_sys_tmp4917 = (r_run_copy8_j_149 + w_sys_intOne);
	assign w_sys_tmp4918 = (r_run_copy9_j_150 + w_sys_intOne);
	assign w_sys_tmp4919 = (r_run_copy10_j_151 + w_sys_intOne);
	assign w_sys_tmp4920 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp5347 = 32'sh00000061;
	assign w_sys_tmp5348 = ( !w_sys_tmp5349 );
	assign w_sys_tmp5349 = (w_sys_tmp5350 < r_run_j_21);
	assign w_sys_tmp5350 = 32'sh00000080;
	assign w_sys_tmp5353 = (w_sys_tmp5354 + w_sys_tmp5356);
	assign w_sys_tmp5354 = (r_run_j_21 * w_sys_tmp5355);
	assign w_sys_tmp5355 = 32'sh00000081;
	assign w_sys_tmp5356 = 32'sh00000021;
	assign w_sys_tmp5357 = w_sub13_result_dataout;
	assign w_sys_tmp5358 = (w_sys_tmp5359 + w_sys_tmp5356);
	assign w_sys_tmp5359 = (r_run_copy10_j_162 * w_sys_tmp5355);
	assign w_sys_tmp5363 = (w_sys_tmp5364 + w_sys_tmp5366);
	assign w_sys_tmp5364 = (r_run_copy9_j_161 * w_sys_tmp5355);
	assign w_sys_tmp5366 = 32'sh00000020;
	assign w_sys_tmp5367 = w_sub12_result_dataout;
	assign w_sys_tmp5368 = (w_sys_tmp5369 + w_sys_tmp5366);
	assign w_sys_tmp5369 = (r_run_copy8_j_160 * w_sys_tmp5355);
	assign w_sys_tmp5373 = (w_sys_tmp5374 + w_sys_tmp5376);
	assign w_sys_tmp5374 = (r_run_copy7_j_159 * w_sys_tmp5355);
	assign w_sys_tmp5376 = 32'sh00000041;
	assign w_sys_tmp5377 = (w_sys_tmp5378 + w_sys_tmp5376);
	assign w_sys_tmp5378 = (r_run_copy6_j_158 * w_sys_tmp5355);
	assign w_sys_tmp5382 = (w_sys_tmp5383 + w_sys_tmp5385);
	assign w_sys_tmp5383 = (r_run_copy5_j_157 * w_sys_tmp5355);
	assign w_sys_tmp5385 = 32'sh00000040;
	assign w_sys_tmp5387 = (w_sys_tmp5388 + w_sys_tmp5385);
	assign w_sys_tmp5388 = (r_run_copy4_j_156 * w_sys_tmp5355);
	assign w_sys_tmp5392 = (w_sys_tmp5393 + w_sys_tmp5395);
	assign w_sys_tmp5393 = (r_run_copy3_j_155 * w_sys_tmp5355);
	assign w_sys_tmp5395 = 32'sh00000061;
	assign w_sys_tmp5396 = (w_sys_tmp5397 + w_sys_tmp5395);
	assign w_sys_tmp5397 = (r_run_copy2_j_154 * w_sys_tmp5355);
	assign w_sys_tmp5401 = (w_sys_tmp5402 + w_sys_tmp5404);
	assign w_sys_tmp5402 = (r_run_copy1_j_153 * w_sys_tmp5355);
	assign w_sys_tmp5404 = 32'sh00000060;
	assign w_sys_tmp5405 = w_sub14_result_dataout;
	assign w_sys_tmp5406 = (w_sys_tmp5407 + w_sys_tmp5404);
	assign w_sys_tmp5407 = (r_run_copy0_j_152 * w_sys_tmp5355);
	assign w_sys_tmp5410 = (r_run_copy0_j_152 + w_sys_intOne);
	assign w_sys_tmp5411 = (r_run_copy1_j_153 + w_sys_intOne);
	assign w_sys_tmp5412 = (r_run_copy2_j_154 + w_sys_intOne);
	assign w_sys_tmp5413 = (r_run_copy3_j_155 + w_sys_intOne);
	assign w_sys_tmp5414 = (r_run_copy4_j_156 + w_sys_intOne);
	assign w_sys_tmp5415 = (r_run_copy5_j_157 + w_sys_intOne);
	assign w_sys_tmp5416 = (r_run_copy6_j_158 + w_sys_intOne);
	assign w_sys_tmp5417 = (r_run_copy7_j_159 + w_sys_intOne);
	assign w_sys_tmp5418 = (r_run_copy8_j_160 + w_sys_intOne);
	assign w_sys_tmp5419 = (r_run_copy9_j_161 + w_sys_intOne);
	assign w_sys_tmp5420 = (r_run_copy10_j_162 + w_sys_intOne);
	assign w_sys_tmp5421 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp5848 = 32'sh00000002;
	assign w_sys_tmp5849 = ( !w_sys_tmp5850 );
	assign w_sys_tmp5850 = (w_sys_tmp5851 < r_run_k_20);
	assign w_sys_tmp5851 = 32'sh00000020;
	assign w_sys_tmp5852 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp5853 = 32'sh00000002;
	assign w_sys_tmp5854 = ( !w_sys_tmp5855 );
	assign w_sys_tmp5855 = (w_sys_tmp5856 < r_run_j_21);
	assign w_sys_tmp5856 = 32'sh00000020;
	assign w_sys_tmp5859 = (w_sys_tmp5860 + r_run_k_20);
	assign w_sys_tmp5860 = (r_run_j_21 * w_sys_tmp5861);
	assign w_sys_tmp5861 = 32'sh00000081;
	assign w_sys_tmp5862 = w_sub00_result_dataout;
	assign w_sys_tmp5863 = (w_sys_tmp5864 + r_run_k_20);
	assign w_sys_tmp5864 = (r_run_copy0_j_163 * w_sys_tmp5861);
	assign w_sys_tmp5866 = (r_run_copy0_j_163 + w_sys_intOne);
	assign w_sys_tmp5867 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp5928 = 32'sh00000021;
	assign w_sys_tmp5929 = ( !w_sys_tmp5930 );
	assign w_sys_tmp5930 = (w_sys_tmp5931 < r_run_j_21);
	assign w_sys_tmp5931 = 32'sh00000040;
	assign w_sys_tmp5934 = (w_sys_tmp5935 + r_run_k_20);
	assign w_sys_tmp5935 = (r_run_j_21 * w_sys_tmp5936);
	assign w_sys_tmp5936 = 32'sh00000081;
	assign w_sys_tmp5937 = w_sub01_result_dataout;
	assign w_sys_tmp5938 = (w_sys_tmp5939 + r_run_k_20);
	assign w_sys_tmp5939 = (r_run_copy0_j_164 * w_sys_tmp5936);
	assign w_sys_tmp5941 = (r_run_copy0_j_164 + w_sys_intOne);
	assign w_sys_tmp5942 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6003 = 32'sh00000041;
	assign w_sys_tmp6004 = ( !w_sys_tmp6005 );
	assign w_sys_tmp6005 = (w_sys_tmp6006 < r_run_j_21);
	assign w_sys_tmp6006 = 32'sh00000060;
	assign w_sys_tmp6009 = (w_sys_tmp6010 + r_run_k_20);
	assign w_sys_tmp6010 = (r_run_j_21 * w_sys_tmp6011);
	assign w_sys_tmp6011 = 32'sh00000081;
	assign w_sys_tmp6012 = w_sub02_result_dataout;
	assign w_sys_tmp6013 = (w_sys_tmp6014 + r_run_k_20);
	assign w_sys_tmp6014 = (r_run_copy0_j_165 * w_sys_tmp6011);
	assign w_sys_tmp6016 = (r_run_copy0_j_165 + w_sys_intOne);
	assign w_sys_tmp6017 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6078 = 32'sh00000061;
	assign w_sys_tmp6079 = ( !w_sys_tmp6080 );
	assign w_sys_tmp6080 = (w_sys_tmp6081 < r_run_j_21);
	assign w_sys_tmp6081 = 32'sh00000080;
	assign w_sys_tmp6084 = (w_sys_tmp6085 + r_run_k_20);
	assign w_sys_tmp6085 = (r_run_j_21 * w_sys_tmp6086);
	assign w_sys_tmp6086 = 32'sh00000081;
	assign w_sys_tmp6087 = w_sub03_result_dataout;
	assign w_sys_tmp6088 = (w_sys_tmp6089 + r_run_k_20);
	assign w_sys_tmp6089 = (r_run_copy0_j_166 * w_sys_tmp6086);
	assign w_sys_tmp6091 = (r_run_copy0_j_166 + w_sys_intOne);
	assign w_sys_tmp6092 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6153 = 32'sh00000021;
	assign w_sys_tmp6154 = ( !w_sys_tmp6155 );
	assign w_sys_tmp6155 = (w_sys_tmp6156 < r_run_k_20);
	assign w_sys_tmp6156 = 32'sh00000040;
	assign w_sys_tmp6157 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp6158 = 32'sh00000002;
	assign w_sys_tmp6159 = ( !w_sys_tmp6160 );
	assign w_sys_tmp6160 = (w_sys_tmp6161 < r_run_j_21);
	assign w_sys_tmp6161 = 32'sh00000020;
	assign w_sys_tmp6164 = (w_sys_tmp6165 + r_run_k_20);
	assign w_sys_tmp6165 = (r_run_j_21 * w_sys_tmp6166);
	assign w_sys_tmp6166 = 32'sh00000081;
	assign w_sys_tmp6167 = w_sub04_result_dataout;
	assign w_sys_tmp6168 = (w_sys_tmp6169 + r_run_k_20);
	assign w_sys_tmp6169 = (r_run_copy0_j_167 * w_sys_tmp6166);
	assign w_sys_tmp6171 = (r_run_copy0_j_167 + w_sys_intOne);
	assign w_sys_tmp6172 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6233 = 32'sh00000021;
	assign w_sys_tmp6234 = ( !w_sys_tmp6235 );
	assign w_sys_tmp6235 = (w_sys_tmp6236 < r_run_j_21);
	assign w_sys_tmp6236 = 32'sh00000040;
	assign w_sys_tmp6239 = (w_sys_tmp6240 + r_run_k_20);
	assign w_sys_tmp6240 = (r_run_j_21 * w_sys_tmp6241);
	assign w_sys_tmp6241 = 32'sh00000081;
	assign w_sys_tmp6242 = w_sub05_result_dataout;
	assign w_sys_tmp6243 = (w_sys_tmp6244 + r_run_k_20);
	assign w_sys_tmp6244 = (r_run_copy0_j_168 * w_sys_tmp6241);
	assign w_sys_tmp6246 = (r_run_copy0_j_168 + w_sys_intOne);
	assign w_sys_tmp6247 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6308 = 32'sh00000041;
	assign w_sys_tmp6309 = ( !w_sys_tmp6310 );
	assign w_sys_tmp6310 = (w_sys_tmp6311 < r_run_j_21);
	assign w_sys_tmp6311 = 32'sh00000060;
	assign w_sys_tmp6314 = (w_sys_tmp6315 + r_run_k_20);
	assign w_sys_tmp6315 = (r_run_j_21 * w_sys_tmp6316);
	assign w_sys_tmp6316 = 32'sh00000081;
	assign w_sys_tmp6317 = w_sub06_result_dataout;
	assign w_sys_tmp6318 = (w_sys_tmp6319 + r_run_k_20);
	assign w_sys_tmp6319 = (r_run_copy0_j_169 * w_sys_tmp6316);
	assign w_sys_tmp6321 = (r_run_copy0_j_169 + w_sys_intOne);
	assign w_sys_tmp6322 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6383 = 32'sh00000061;
	assign w_sys_tmp6384 = ( !w_sys_tmp6385 );
	assign w_sys_tmp6385 = (w_sys_tmp6386 < r_run_j_21);
	assign w_sys_tmp6386 = 32'sh00000080;
	assign w_sys_tmp6389 = (w_sys_tmp6390 + r_run_k_20);
	assign w_sys_tmp6390 = (r_run_j_21 * w_sys_tmp6391);
	assign w_sys_tmp6391 = 32'sh00000081;
	assign w_sys_tmp6392 = w_sub07_result_dataout;
	assign w_sys_tmp6393 = (w_sys_tmp6394 + r_run_k_20);
	assign w_sys_tmp6394 = (r_run_copy0_j_170 * w_sys_tmp6391);
	assign w_sys_tmp6396 = (r_run_copy0_j_170 + w_sys_intOne);
	assign w_sys_tmp6397 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6458 = 32'sh00000041;
	assign w_sys_tmp6459 = ( !w_sys_tmp6460 );
	assign w_sys_tmp6460 = (w_sys_tmp6461 < r_run_k_20);
	assign w_sys_tmp6461 = 32'sh00000060;
	assign w_sys_tmp6462 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp6463 = 32'sh00000002;
	assign w_sys_tmp6464 = ( !w_sys_tmp6465 );
	assign w_sys_tmp6465 = (w_sys_tmp6466 < r_run_j_21);
	assign w_sys_tmp6466 = 32'sh00000020;
	assign w_sys_tmp6469 = (w_sys_tmp6470 + r_run_k_20);
	assign w_sys_tmp6470 = (r_run_j_21 * w_sys_tmp6471);
	assign w_sys_tmp6471 = 32'sh00000081;
	assign w_sys_tmp6472 = w_sub08_result_dataout;
	assign w_sys_tmp6473 = (w_sys_tmp6474 + r_run_k_20);
	assign w_sys_tmp6474 = (r_run_copy0_j_171 * w_sys_tmp6471);
	assign w_sys_tmp6476 = (r_run_copy0_j_171 + w_sys_intOne);
	assign w_sys_tmp6477 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6538 = 32'sh00000021;
	assign w_sys_tmp6539 = ( !w_sys_tmp6540 );
	assign w_sys_tmp6540 = (w_sys_tmp6541 < r_run_j_21);
	assign w_sys_tmp6541 = 32'sh00000040;
	assign w_sys_tmp6544 = (w_sys_tmp6545 + r_run_k_20);
	assign w_sys_tmp6545 = (r_run_j_21 * w_sys_tmp6546);
	assign w_sys_tmp6546 = 32'sh00000081;
	assign w_sys_tmp6547 = w_sub09_result_dataout;
	assign w_sys_tmp6548 = (w_sys_tmp6549 + r_run_k_20);
	assign w_sys_tmp6549 = (r_run_copy0_j_172 * w_sys_tmp6546);
	assign w_sys_tmp6551 = (r_run_copy0_j_172 + w_sys_intOne);
	assign w_sys_tmp6552 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6613 = 32'sh00000041;
	assign w_sys_tmp6614 = ( !w_sys_tmp6615 );
	assign w_sys_tmp6615 = (w_sys_tmp6616 < r_run_j_21);
	assign w_sys_tmp6616 = 32'sh00000060;
	assign w_sys_tmp6619 = (w_sys_tmp6620 + r_run_k_20);
	assign w_sys_tmp6620 = (r_run_j_21 * w_sys_tmp6621);
	assign w_sys_tmp6621 = 32'sh00000081;
	assign w_sys_tmp6622 = w_sub10_result_dataout;
	assign w_sys_tmp6623 = (w_sys_tmp6624 + r_run_k_20);
	assign w_sys_tmp6624 = (r_run_copy0_j_173 * w_sys_tmp6621);
	assign w_sys_tmp6626 = (r_run_copy0_j_173 + w_sys_intOne);
	assign w_sys_tmp6627 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6688 = 32'sh00000061;
	assign w_sys_tmp6689 = ( !w_sys_tmp6690 );
	assign w_sys_tmp6690 = (w_sys_tmp6691 < r_run_j_21);
	assign w_sys_tmp6691 = 32'sh00000080;
	assign w_sys_tmp6694 = (w_sys_tmp6695 + r_run_k_20);
	assign w_sys_tmp6695 = (r_run_j_21 * w_sys_tmp6696);
	assign w_sys_tmp6696 = 32'sh00000081;
	assign w_sys_tmp6697 = w_sub11_result_dataout;
	assign w_sys_tmp6698 = (w_sys_tmp6699 + r_run_k_20);
	assign w_sys_tmp6699 = (r_run_copy0_j_174 * w_sys_tmp6696);
	assign w_sys_tmp6701 = (r_run_copy0_j_174 + w_sys_intOne);
	assign w_sys_tmp6702 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6763 = 32'sh00000061;
	assign w_sys_tmp6764 = ( !w_sys_tmp6765 );
	assign w_sys_tmp6765 = (w_sys_tmp6766 < r_run_k_20);
	assign w_sys_tmp6766 = 32'sh00000080;
	assign w_sys_tmp6767 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp6768 = 32'sh00000002;
	assign w_sys_tmp6769 = ( !w_sys_tmp6770 );
	assign w_sys_tmp6770 = (w_sys_tmp6771 < r_run_j_21);
	assign w_sys_tmp6771 = 32'sh00000020;
	assign w_sys_tmp6774 = (w_sys_tmp6775 + r_run_k_20);
	assign w_sys_tmp6775 = (r_run_j_21 * w_sys_tmp6776);
	assign w_sys_tmp6776 = 32'sh00000081;
	assign w_sys_tmp6777 = w_sub12_result_dataout;
	assign w_sys_tmp6778 = (w_sys_tmp6779 + r_run_k_20);
	assign w_sys_tmp6779 = (r_run_copy0_j_175 * w_sys_tmp6776);
	assign w_sys_tmp6781 = (r_run_copy0_j_175 + w_sys_intOne);
	assign w_sys_tmp6782 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6843 = 32'sh00000021;
	assign w_sys_tmp6844 = ( !w_sys_tmp6845 );
	assign w_sys_tmp6845 = (w_sys_tmp6846 < r_run_j_21);
	assign w_sys_tmp6846 = 32'sh00000040;
	assign w_sys_tmp6849 = (w_sys_tmp6850 + r_run_k_20);
	assign w_sys_tmp6850 = (r_run_j_21 * w_sys_tmp6851);
	assign w_sys_tmp6851 = 32'sh00000081;
	assign w_sys_tmp6852 = w_sub13_result_dataout;
	assign w_sys_tmp6853 = (w_sys_tmp6854 + r_run_k_20);
	assign w_sys_tmp6854 = (r_run_copy0_j_176 * w_sys_tmp6851);
	assign w_sys_tmp6856 = (r_run_copy0_j_176 + w_sys_intOne);
	assign w_sys_tmp6857 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6918 = 32'sh00000041;
	assign w_sys_tmp6919 = ( !w_sys_tmp6920 );
	assign w_sys_tmp6920 = (w_sys_tmp6921 < r_run_j_21);
	assign w_sys_tmp6921 = 32'sh00000060;
	assign w_sys_tmp6924 = (w_sys_tmp6925 + r_run_k_20);
	assign w_sys_tmp6925 = (r_run_j_21 * w_sys_tmp6926);
	assign w_sys_tmp6926 = 32'sh00000081;
	assign w_sys_tmp6927 = w_sub14_result_dataout;
	assign w_sys_tmp6928 = (w_sys_tmp6929 + r_run_k_20);
	assign w_sys_tmp6929 = (r_run_copy0_j_177 * w_sys_tmp6926);
	assign w_sys_tmp6931 = (r_run_copy0_j_177 + w_sys_intOne);
	assign w_sys_tmp6932 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6993 = 32'sh00000061;
	assign w_sys_tmp6994 = ( !w_sys_tmp6995 );
	assign w_sys_tmp6995 = (w_sys_tmp6996 < r_run_j_21);
	assign w_sys_tmp6996 = 32'sh00000080;
	assign w_sys_tmp6999 = (w_sys_tmp7000 + r_run_k_20);
	assign w_sys_tmp7000 = (r_run_j_21 * w_sys_tmp7001);
	assign w_sys_tmp7001 = 32'sh00000081;
	assign w_sys_tmp7002 = w_sub15_result_dataout;
	assign w_sys_tmp7003 = (w_sys_tmp7004 + r_run_k_20);
	assign w_sys_tmp7004 = (r_run_copy0_j_178 * w_sys_tmp7001);
	assign w_sys_tmp7006 = (r_run_copy0_j_178 + w_sys_intOne);
	assign w_sys_tmp7007 = (r_run_j_21 + w_sys_intOne);


	sub09
		sub09_inst(
			.i_fld_T_0_addr_0 (w_sub09_T_addr),
			.i_fld_T_0_datain_0 (w_sub09_T_datain),
			.o_fld_T_0_dataout_0 (w_sub09_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub09_T_r_w),
			.i_fld_U_2_addr_0 (w_sub09_U_addr),
			.i_fld_U_2_datain_0 (w_sub09_U_datain),
			.o_fld_U_2_dataout_0 (w_sub09_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub09_U_r_w),
			.i_fld_V_1_addr_0 (w_sub09_V_addr),
			.i_fld_V_1_datain_0 (w_sub09_V_datain),
			.o_fld_V_1_dataout_0 (w_sub09_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub09_V_r_w),
			.i_fld_result_3_addr_0 (w_sub09_result_addr),
			.i_fld_result_3_datain_0 (w_sub09_result_datain),
			.o_fld_result_3_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub09_result_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_T_0_addr_0 (w_sub08_T_addr),
			.i_fld_T_0_datain_0 (w_sub08_T_datain),
			.o_fld_T_0_dataout_0 (w_sub08_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub08_T_r_w),
			.i_fld_U_2_addr_0 (w_sub08_U_addr),
			.i_fld_U_2_datain_0 (w_sub08_U_datain),
			.o_fld_U_2_dataout_0 (w_sub08_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub08_U_r_w),
			.i_fld_V_1_addr_0 (w_sub08_V_addr),
			.i_fld_V_1_datain_0 (w_sub08_V_datain),
			.o_fld_V_1_dataout_0 (w_sub08_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub08_V_r_w),
			.i_fld_result_3_addr_0 (w_sub08_result_addr),
			.i_fld_result_3_datain_0 (w_sub08_result_datain),
			.o_fld_result_3_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub08_result_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_T_0_addr_0 (w_sub12_T_addr),
			.i_fld_T_0_datain_0 (w_sub12_T_datain),
			.o_fld_T_0_dataout_0 (w_sub12_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub12_T_r_w),
			.i_fld_U_2_addr_0 (w_sub12_U_addr),
			.i_fld_U_2_datain_0 (w_sub12_U_datain),
			.o_fld_U_2_dataout_0 (w_sub12_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub12_U_r_w),
			.i_fld_V_1_addr_0 (w_sub12_V_addr),
			.i_fld_V_1_datain_0 (w_sub12_V_datain),
			.o_fld_V_1_dataout_0 (w_sub12_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub12_V_r_w),
			.i_fld_result_3_addr_0 (w_sub12_result_addr),
			.i_fld_result_3_datain_0 (w_sub12_result_datain),
			.o_fld_result_3_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub12_result_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_T_0_addr_0 (w_sub03_T_addr),
			.i_fld_T_0_datain_0 (w_sub03_T_datain),
			.o_fld_T_0_dataout_0 (w_sub03_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub03_T_r_w),
			.i_fld_U_2_addr_0 (w_sub03_U_addr),
			.i_fld_U_2_datain_0 (w_sub03_U_datain),
			.o_fld_U_2_dataout_0 (w_sub03_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub03_U_r_w),
			.i_fld_V_1_addr_0 (w_sub03_V_addr),
			.i_fld_V_1_datain_0 (w_sub03_V_datain),
			.o_fld_V_1_dataout_0 (w_sub03_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub03_V_r_w),
			.i_fld_result_3_addr_0 (w_sub03_result_addr),
			.i_fld_result_3_datain_0 (w_sub03_result_datain),
			.o_fld_result_3_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub03_result_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_T_0_addr_0 (w_sub02_T_addr),
			.i_fld_T_0_datain_0 (w_sub02_T_datain),
			.o_fld_T_0_dataout_0 (w_sub02_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub02_T_r_w),
			.i_fld_U_2_addr_0 (w_sub02_U_addr),
			.i_fld_U_2_datain_0 (w_sub02_U_datain),
			.o_fld_U_2_dataout_0 (w_sub02_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub02_U_r_w),
			.i_fld_V_1_addr_0 (w_sub02_V_addr),
			.i_fld_V_1_datain_0 (w_sub02_V_datain),
			.o_fld_V_1_dataout_0 (w_sub02_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub02_V_r_w),
			.i_fld_result_3_addr_0 (w_sub02_result_addr),
			.i_fld_result_3_datain_0 (w_sub02_result_datain),
			.o_fld_result_3_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub02_result_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_T_0_addr_0 (w_sub11_T_addr),
			.i_fld_T_0_datain_0 (w_sub11_T_datain),
			.o_fld_T_0_dataout_0 (w_sub11_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub11_T_r_w),
			.i_fld_U_2_addr_0 (w_sub11_U_addr),
			.i_fld_U_2_datain_0 (w_sub11_U_datain),
			.o_fld_U_2_dataout_0 (w_sub11_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub11_U_r_w),
			.i_fld_V_1_addr_0 (w_sub11_V_addr),
			.i_fld_V_1_datain_0 (w_sub11_V_datain),
			.o_fld_V_1_dataout_0 (w_sub11_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub11_V_r_w),
			.i_fld_result_3_addr_0 (w_sub11_result_addr),
			.i_fld_result_3_datain_0 (w_sub11_result_datain),
			.o_fld_result_3_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub11_result_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_T_0_addr_0 (w_sub14_T_addr),
			.i_fld_T_0_datain_0 (w_sub14_T_datain),
			.o_fld_T_0_dataout_0 (w_sub14_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub14_T_r_w),
			.i_fld_U_2_addr_0 (w_sub14_U_addr),
			.i_fld_U_2_datain_0 (w_sub14_U_datain),
			.o_fld_U_2_dataout_0 (w_sub14_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub14_U_r_w),
			.i_fld_V_1_addr_0 (w_sub14_V_addr),
			.i_fld_V_1_datain_0 (w_sub14_V_datain),
			.o_fld_V_1_dataout_0 (w_sub14_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub14_V_r_w),
			.i_fld_result_3_addr_0 (w_sub14_result_addr),
			.i_fld_result_3_datain_0 (w_sub14_result_datain),
			.o_fld_result_3_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub14_result_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_T_0_addr_0 (w_sub01_T_addr),
			.i_fld_T_0_datain_0 (w_sub01_T_datain),
			.o_fld_T_0_dataout_0 (w_sub01_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub01_T_r_w),
			.i_fld_U_2_addr_0 (w_sub01_U_addr),
			.i_fld_U_2_datain_0 (w_sub01_U_datain),
			.o_fld_U_2_dataout_0 (w_sub01_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub01_U_r_w),
			.i_fld_V_1_addr_0 (w_sub01_V_addr),
			.i_fld_V_1_datain_0 (w_sub01_V_datain),
			.o_fld_V_1_dataout_0 (w_sub01_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub01_V_r_w),
			.i_fld_result_3_addr_0 (w_sub01_result_addr),
			.i_fld_result_3_datain_0 (w_sub01_result_datain),
			.o_fld_result_3_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub01_result_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_T_0_addr_0 (w_sub13_T_addr),
			.i_fld_T_0_datain_0 (w_sub13_T_datain),
			.o_fld_T_0_dataout_0 (w_sub13_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub13_T_r_w),
			.i_fld_U_2_addr_0 (w_sub13_U_addr),
			.i_fld_U_2_datain_0 (w_sub13_U_datain),
			.o_fld_U_2_dataout_0 (w_sub13_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub13_U_r_w),
			.i_fld_V_1_addr_0 (w_sub13_V_addr),
			.i_fld_V_1_datain_0 (w_sub13_V_datain),
			.o_fld_V_1_dataout_0 (w_sub13_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub13_V_r_w),
			.i_fld_result_3_addr_0 (w_sub13_result_addr),
			.i_fld_result_3_datain_0 (w_sub13_result_datain),
			.o_fld_result_3_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub13_result_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_T_0_addr_0 (w_sub00_T_addr),
			.i_fld_T_0_datain_0 (w_sub00_T_datain),
			.o_fld_T_0_dataout_0 (w_sub00_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub00_T_r_w),
			.i_fld_U_2_addr_0 (w_sub00_U_addr),
			.i_fld_U_2_datain_0 (w_sub00_U_datain),
			.o_fld_U_2_dataout_0 (w_sub00_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub00_U_r_w),
			.i_fld_V_1_addr_0 (w_sub00_V_addr),
			.i_fld_V_1_datain_0 (w_sub00_V_datain),
			.o_fld_V_1_dataout_0 (w_sub00_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub00_V_r_w),
			.i_fld_result_3_addr_0 (w_sub00_result_addr),
			.i_fld_result_3_datain_0 (w_sub00_result_datain),
			.o_fld_result_3_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub00_result_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_T_0_addr_0 (w_sub07_T_addr),
			.i_fld_T_0_datain_0 (w_sub07_T_datain),
			.o_fld_T_0_dataout_0 (w_sub07_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub07_T_r_w),
			.i_fld_U_2_addr_0 (w_sub07_U_addr),
			.i_fld_U_2_datain_0 (w_sub07_U_datain),
			.o_fld_U_2_dataout_0 (w_sub07_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub07_U_r_w),
			.i_fld_V_1_addr_0 (w_sub07_V_addr),
			.i_fld_V_1_datain_0 (w_sub07_V_datain),
			.o_fld_V_1_dataout_0 (w_sub07_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub07_V_r_w),
			.i_fld_result_3_addr_0 (w_sub07_result_addr),
			.i_fld_result_3_datain_0 (w_sub07_result_datain),
			.o_fld_result_3_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub07_result_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_T_0_addr_0 (w_sub06_T_addr),
			.i_fld_T_0_datain_0 (w_sub06_T_datain),
			.o_fld_T_0_dataout_0 (w_sub06_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub06_T_r_w),
			.i_fld_U_2_addr_0 (w_sub06_U_addr),
			.i_fld_U_2_datain_0 (w_sub06_U_datain),
			.o_fld_U_2_dataout_0 (w_sub06_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub06_U_r_w),
			.i_fld_V_1_addr_0 (w_sub06_V_addr),
			.i_fld_V_1_datain_0 (w_sub06_V_datain),
			.o_fld_V_1_dataout_0 (w_sub06_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub06_V_r_w),
			.i_fld_result_3_addr_0 (w_sub06_result_addr),
			.i_fld_result_3_datain_0 (w_sub06_result_datain),
			.o_fld_result_3_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub06_result_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_T_0_addr_0 (w_sub15_T_addr),
			.i_fld_T_0_datain_0 (w_sub15_T_datain),
			.o_fld_T_0_dataout_0 (w_sub15_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub15_T_r_w),
			.i_fld_U_2_addr_0 (w_sub15_U_addr),
			.i_fld_U_2_datain_0 (w_sub15_U_datain),
			.o_fld_U_2_dataout_0 (w_sub15_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub15_U_r_w),
			.i_fld_V_1_addr_0 (w_sub15_V_addr),
			.i_fld_V_1_datain_0 (w_sub15_V_datain),
			.o_fld_V_1_dataout_0 (w_sub15_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub15_V_r_w),
			.i_fld_result_3_addr_0 (w_sub15_result_addr),
			.i_fld_result_3_datain_0 (w_sub15_result_datain),
			.o_fld_result_3_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub15_result_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_T_0_addr_0 (w_sub05_T_addr),
			.i_fld_T_0_datain_0 (w_sub05_T_datain),
			.o_fld_T_0_dataout_0 (w_sub05_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub05_T_r_w),
			.i_fld_U_2_addr_0 (w_sub05_U_addr),
			.i_fld_U_2_datain_0 (w_sub05_U_datain),
			.o_fld_U_2_dataout_0 (w_sub05_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub05_U_r_w),
			.i_fld_V_1_addr_0 (w_sub05_V_addr),
			.i_fld_V_1_datain_0 (w_sub05_V_datain),
			.o_fld_V_1_dataout_0 (w_sub05_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub05_V_r_w),
			.i_fld_result_3_addr_0 (w_sub05_result_addr),
			.i_fld_result_3_datain_0 (w_sub05_result_datain),
			.o_fld_result_3_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub05_result_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_T_0_addr_0 (w_sub04_T_addr),
			.i_fld_T_0_datain_0 (w_sub04_T_datain),
			.o_fld_T_0_dataout_0 (w_sub04_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub04_T_r_w),
			.i_fld_U_2_addr_0 (w_sub04_U_addr),
			.i_fld_U_2_datain_0 (w_sub04_U_datain),
			.o_fld_U_2_dataout_0 (w_sub04_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub04_U_r_w),
			.i_fld_V_1_addr_0 (w_sub04_V_addr),
			.i_fld_V_1_datain_0 (w_sub04_V_datain),
			.o_fld_V_1_dataout_0 (w_sub04_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub04_V_r_w),
			.i_fld_result_3_addr_0 (w_sub04_result_addr),
			.i_fld_result_3_datain_0 (w_sub04_result_datain),
			.o_fld_result_3_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub04_result_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_T_0_addr_0 (w_sub10_T_addr),
			.i_fld_T_0_datain_0 (w_sub10_T_datain),
			.o_fld_T_0_dataout_0 (w_sub10_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub10_T_r_w),
			.i_fld_U_2_addr_0 (w_sub10_U_addr),
			.i_fld_U_2_datain_0 (w_sub10_U_datain),
			.o_fld_U_2_dataout_0 (w_sub10_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub10_U_r_w),
			.i_fld_V_1_addr_0 (w_sub10_V_addr),
			.i_fld_V_1_datain_0 (w_sub10_V_datain),
			.o_fld_V_1_dataout_0 (w_sub10_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub10_V_r_w),
			.i_fld_result_3_addr_0 (w_sub10_result_addr),
			.i_fld_result_3_datain_0 (w_sub10_result_datain),
			.o_fld_result_3_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub10_result_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_V_3(
			.clk (clock),
			.ce_0 (w_fld_V_3_ce_0),
			.addr_0 (w_fld_V_3_addr_0),
			.datain_0 (w_fld_V_3_datain_0),
			.dataout_0 (w_fld_V_3_dataout_0),
			.r_w_0 (w_fld_V_3_r_w_0),
			.ce_1 (w_fld_V_3_ce_1),
			.addr_1 (r_fld_V_3_addr_1),
			.datain_1 (r_fld_V_3_datain_1),
			.dataout_1 (w_fld_V_3_dataout_1),
			.r_w_1 (r_fld_V_3_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp38;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==6'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h18)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h16)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp36;

									end
									else
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp18;

									end
									else
									if((6'h7<=r_sys_run_step && r_sys_run_step<=6'hb) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'hf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_27;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h7<=r_sys_run_step && r_sys_run_step<=6'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h16)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_32;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp37;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						9'h12f: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 9'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h0: begin
							r_sys_run_phase <= 9'h2;
						end

						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h4;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h5;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12) ? 9'h9 : 9'hf);

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h5;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'ha;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp15) ? 9'hd : 9'h6);

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_phase <= 9'ha;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h10;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp226) ? 9'h14 : 9'h2c);

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h10;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h15;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp230) ? 9'h18 : 9'h1a);

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h15;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h1b;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp445) ? 9'h1e : 9'h20);

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h1b;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h21;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp660) ? 9'h24 : 9'h26);

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h21;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h27;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp875) ? 9'h2a : 9'h11);

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h27;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h2d;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1090) ? 9'h31 : 9'h49);

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h2d;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h32;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1094) ? 9'h35 : 9'h37);

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h32;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h38;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1309) ? 9'h3b : 9'h3d);

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h38;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h3e;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1524) ? 9'h41 : 9'h43);

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h3e;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h44;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1739) ? 9'h47 : 9'h2e);

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h44;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h4a;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1954) ? 9'h4e : 9'h66);

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h4a;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h4f;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1958) ? 9'h52 : 9'h54);

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h4f;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h55;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2173) ? 9'h58 : 9'h5a);

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h55;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h5b;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2388) ? 9'h5e : 9'h60);

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h5b;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h61;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2603) ? 9'h64 : 9'h4b);

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h61;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h67;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2818) ? 9'h6b : 9'h83);

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h67;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h6c;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2822) ? 9'h6f : 9'h71);

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h6c;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h72;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3037) ? 9'h75 : 9'h77);

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h72;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h78;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3252) ? 9'h7b : 9'h7d);

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h78;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h7e;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3467) ? 9'h81 : 9'h68);

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h7e;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h84;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3681) ? 9'h87 : 9'hbb);

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h84;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 9'h89;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 9'h8b;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h8c;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3685) ? 9'h8f : 9'h91);

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_phase <= 9'h8c;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h92;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3725) ? 9'h95 : 9'h97);

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_phase <= 9'h92;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h98;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3765) ? 9'h9b : 9'h9d);

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_phase <= 9'h98;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h9e;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3805) ? 9'ha1 : 9'ha3);

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_phase <= 9'h9e;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'ha4;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3845) ? 9'ha7 : 9'ha9);

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 9'ha4;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'haa;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4346) ? 9'had : 9'haf);

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 9'haa;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hb0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4847) ? 9'hb3 : 9'hb5);

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 9'hb0;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hb6;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5348) ? 9'hb9 : 9'h85);

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 9'hb6;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hbc;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5849) ? 9'hc0 : 9'hd8);

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hbc;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hc1;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5854) ? 9'hc4 : 9'hc6);

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hc1;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hc7;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5929) ? 9'hca : 9'hcc);

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hc7;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hcd;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6004) ? 9'hd0 : 9'hd2);

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hcd;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hd3;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6079) ? 9'hd6 : 9'hbd);

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hd3;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hd9;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6154) ? 9'hdd : 9'hf5);

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hd9;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hde;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6159) ? 9'he1 : 9'he3);

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hde;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'he4;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6234) ? 9'he7 : 9'he9);

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'he4;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hea;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6309) ? 9'hed : 9'hef);

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hea;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hf0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6384) ? 9'hf3 : 9'hda);

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hf0;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hf6;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6459) ? 9'hfa : 9'h112);

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hf6;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'hfb;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6464) ? 9'hfe : 9'h100);

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'hfb;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h101;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6539) ? 9'h104 : 9'h106);

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h101;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h107;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6614) ? 9'h10a : 9'h10c);

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h107;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h10d;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6689) ? 9'h110 : 9'hf7);

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h10d;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h113;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6764) ? 9'h117 : 9'h12f);

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h113;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h118;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6769) ? 9'h11b : 9'h11d);

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h118;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h11e;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6844) ? 9'h121 : 9'h123);

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h11e;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h124;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6919) ? 9'h127 : 9'h129);

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h124;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 9'h12a;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6994) ? 9'h12d : 9'h114);

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 9'h12a;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sys_run_phase <= 9'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						9'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						9'h12f: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp22[14:0] );

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp255[14:0] );

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp470[14:0] );

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp685[14:0] );

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp900[14:0] );

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1119[14:0] );

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1334[14:0] );

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1549[14:0] );

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1764[14:0] );

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1983[14:0] );

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2198[14:0] );

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2413[14:0] );

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2628[14:0] );

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2847[14:0] );

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3062[14:0] );

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3277[14:0] );

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3492[14:0] );

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp5859[14:0] );

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp5934[14:0] );

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6009[14:0] );

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6084[14:0] );

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6164[14:0] );

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6239[14:0] );

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6314[14:0] );

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6389[14:0] );

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6469[14:0] );

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6544[14:0] );

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6619[14:0] );

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6694[14:0] );

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6774[14:0] );

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6849[14:0] );

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6924[14:0] );

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6999[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp5862;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp5937;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6012;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6087;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6167;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6242;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6317;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6392;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6472;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6547;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6622;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6697;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6777;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6852;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6927;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp7002;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12f: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp27[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12f: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp32[14:0] );

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp239[14:0] );

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp454[14:0] );

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp669[14:0] );

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp884[14:0] );

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1103[14:0] );

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1318[14:0] );

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1533[14:0] );

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1748[14:0] );

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1967[14:0] );

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2182[14:0] );

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2397[14:0] );

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2612[14:0] );

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2831[14:0] );

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3046[14:0] );

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3261[14:0] );

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3476[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp41[14:0] );

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp247[14:0] );

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp462[14:0] );

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp677[14:0] );

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp892[14:0] );

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1111[14:0] );

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1326[14:0] );

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1541[14:0] );

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1756[14:0] );

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1975[14:0] );

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2190[14:0] );

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2405[14:0] );

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2620[14:0] );

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2839[14:0] );

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3054[14:0] );

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3269[14:0] );

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3484[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_fld_V_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp14;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp229;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp1089;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp1093;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp1953;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp1957;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp2817;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp2821;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp3684;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_run_k_20 <= w_sys_tmp3723;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp3724;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_run_k_20 <= w_sys_tmp3763;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp3764;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_run_k_20 <= w_sys_tmp3803;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp3804;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_run_k_20 <= w_sys_tmp3843;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp5848;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp5852;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp6153;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp6157;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp6458;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp6462;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp6763;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_20 <= w_sys_tmp6767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_21 <= w_sys_tmp48;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp263;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp444;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp478;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp659;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp693;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp874;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp908;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp1127;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp1308;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp1342;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp1523;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp1557;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp1738;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp1772;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp1991;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp2172;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp2206;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp2387;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp2421;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp2602;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp2636;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp2855;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp3036;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp3070;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp3251;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp3285;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp3466;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp3500;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp3844;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_21 <= w_sys_tmp3918;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp4345;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_21 <= w_sys_tmp4419;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp4846;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_21 <= w_sys_tmp4920;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp5347;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_21 <= w_sys_tmp5421;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp5853;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp5867;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp5928;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp5942;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6003;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6017;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6078;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6092;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6158;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6172;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6233;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6247;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6308;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6322;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6383;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6397;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6463;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6477;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6538;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6552;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6613;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6627;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6688;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6702;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6768;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6782;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6843;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6857;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6918;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp6932;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_21 <= w_sys_tmp6993;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_21 <= w_sys_tmp7007;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_22 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_22 <= w_sys_tmp3683;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_mx_23 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_my_24 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dt_25 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dx_26 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dy_27 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r1_28 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r2_29 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r3_30 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r4_31 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h11)) begin
										r_run_YY_32 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14)) begin
										r_run_YY_32 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_kx_33 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_ky_34 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_nlast_35 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_36 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_36 <= w_sys_tmp45;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_37 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_run_copy1_j_37 <= w_sys_tmp46;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_38 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_38 <= w_sys_tmp47;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_39 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_39 <= w_sys_tmp258;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_40 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_40 <= w_sys_tmp259;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_41 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_41 <= w_sys_tmp260;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_42 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_42 <= w_sys_tmp261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_43 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_43 <= w_sys_tmp262;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_44 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_44 <= w_sys_tmp473;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_45 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_45 <= w_sys_tmp474;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_46 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_46 <= w_sys_tmp475;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_47 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_47 <= w_sys_tmp476;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_48 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_48 <= w_sys_tmp477;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_49 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_49 <= w_sys_tmp688;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_50 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_50 <= w_sys_tmp689;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_51 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_51 <= w_sys_tmp690;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_52 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_52 <= w_sys_tmp691;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_53 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_53 <= w_sys_tmp692;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_54 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_54 <= w_sys_tmp903;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_55 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_55 <= w_sys_tmp904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_56 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_56 <= w_sys_tmp905;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_57 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_57 <= w_sys_tmp906;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_58 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_58 <= w_sys_tmp907;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_59 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_59 <= w_sys_tmp1122;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_60 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_60 <= w_sys_tmp1123;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_61 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_61 <= w_sys_tmp1124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_62 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_62 <= w_sys_tmp1125;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_63 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_63 <= w_sys_tmp1126;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_64 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_64 <= w_sys_tmp1337;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_65 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_65 <= w_sys_tmp1338;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_66 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_66 <= w_sys_tmp1339;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_67 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_67 <= w_sys_tmp1340;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_68 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_68 <= w_sys_tmp1341;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_69 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_69 <= w_sys_tmp1552;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_70 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_70 <= w_sys_tmp1553;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_71 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_71 <= w_sys_tmp1554;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_72 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_72 <= w_sys_tmp1555;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_73 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_73 <= w_sys_tmp1556;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_74 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_74 <= w_sys_tmp1767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_75 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_75 <= w_sys_tmp1768;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_76 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_76 <= w_sys_tmp1769;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_77 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_77 <= w_sys_tmp1770;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_78 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_78 <= w_sys_tmp1771;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_79 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_79 <= w_sys_tmp1986;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_80 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_80 <= w_sys_tmp1987;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_81 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_81 <= w_sys_tmp1988;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_82 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_82 <= w_sys_tmp1989;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_83 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_83 <= w_sys_tmp1990;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_84 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_84 <= w_sys_tmp2201;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_85 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_85 <= w_sys_tmp2202;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_86 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_86 <= w_sys_tmp2203;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_87 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_87 <= w_sys_tmp2204;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_88 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_88 <= w_sys_tmp2205;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_89 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_89 <= w_sys_tmp2416;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_90 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_90 <= w_sys_tmp2417;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_91 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_91 <= w_sys_tmp2418;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_92 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_92 <= w_sys_tmp2419;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_93 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_93 <= w_sys_tmp2420;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_94 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_94 <= w_sys_tmp2631;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_95 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_95 <= w_sys_tmp2632;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_96 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_96 <= w_sys_tmp2633;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_97 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_97 <= w_sys_tmp2634;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_98 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_98 <= w_sys_tmp2635;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_99 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_99 <= w_sys_tmp2850;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_100 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_100 <= w_sys_tmp2851;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_101 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_101 <= w_sys_tmp2852;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_102 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_102 <= w_sys_tmp2853;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_103 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_103 <= w_sys_tmp2854;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_104 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_104 <= w_sys_tmp3065;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_105 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_105 <= w_sys_tmp3066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_106 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_106 <= w_sys_tmp3067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_107 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_107 <= w_sys_tmp3068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_108 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_108 <= w_sys_tmp3069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_109 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_109 <= w_sys_tmp3280;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_110 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_110 <= w_sys_tmp3281;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_111 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_111 <= w_sys_tmp3282;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_112 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_112 <= w_sys_tmp3283;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_113 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_113 <= w_sys_tmp3284;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_114 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_114 <= w_sys_tmp3495;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_115 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_115 <= w_sys_tmp3496;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_116 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_116 <= w_sys_tmp3497;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_117 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_117 <= w_sys_tmp3498;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_118 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_118 <= w_sys_tmp3499;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_119 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_119 <= w_sys_tmp3907;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_120 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_120 <= w_sys_tmp3908;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_121 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_121 <= w_sys_tmp3909;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_122 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_122 <= w_sys_tmp3910;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_123 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_123 <= w_sys_tmp3911;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_124 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_124 <= w_sys_tmp3912;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_125 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_125 <= w_sys_tmp3913;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_126 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_126 <= w_sys_tmp3914;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_127 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_127 <= w_sys_tmp3915;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_128 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_128 <= w_sys_tmp3916;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_129 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_129 <= w_sys_tmp3917;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_130 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_130 <= w_sys_tmp4408;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_131 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_131 <= w_sys_tmp4409;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_132 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_132 <= w_sys_tmp4410;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_133 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_133 <= w_sys_tmp4411;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_134 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_134 <= w_sys_tmp4412;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_135 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_135 <= w_sys_tmp4413;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_136 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_136 <= w_sys_tmp4414;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_137 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_137 <= w_sys_tmp4415;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_138 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_138 <= w_sys_tmp4416;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_139 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_139 <= w_sys_tmp4417;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_140 <= r_run_j_21;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_140 <= w_sys_tmp4418;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_141 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_141 <= w_sys_tmp4909;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_142 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_142 <= w_sys_tmp4910;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_143 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_143 <= w_sys_tmp4911;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_144 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_144 <= w_sys_tmp4912;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_145 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_145 <= w_sys_tmp4913;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_146 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_146 <= w_sys_tmp4914;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_147 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_147 <= w_sys_tmp4915;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_148 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_148 <= w_sys_tmp4916;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_149 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_149 <= w_sys_tmp4917;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_150 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_150 <= w_sys_tmp4918;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_151 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_151 <= w_sys_tmp4919;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_152 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_152 <= w_sys_tmp5410;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_153 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_153 <= w_sys_tmp5411;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_154 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_154 <= w_sys_tmp5412;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_155 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_155 <= w_sys_tmp5413;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_156 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_156 <= w_sys_tmp5414;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_157 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_157 <= w_sys_tmp5415;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_158 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_158 <= w_sys_tmp5416;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_159 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_159 <= w_sys_tmp5417;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_160 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_160 <= w_sys_tmp5418;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_161 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_161 <= w_sys_tmp5419;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_162 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_162 <= w_sys_tmp5420;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_163 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_163 <= w_sys_tmp5866;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_164 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_164 <= w_sys_tmp5941;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hcc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_165 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_165 <= w_sys_tmp6016;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_166 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_166 <= w_sys_tmp6091;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_167 <= r_run_j_21;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_167 <= w_sys_tmp6171;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_168 <= r_run_j_21;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_168 <= w_sys_tmp6246;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_169 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_169 <= w_sys_tmp6321;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_170 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_170 <= w_sys_tmp6396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hfa: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_171 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_171 <= w_sys_tmp6476;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h100: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_172 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_172 <= w_sys_tmp6551;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h106: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_173 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_173 <= w_sys_tmp6626;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h10c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_174 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_174 <= w_sys_tmp6701;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h117: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_175 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_175 <= w_sys_tmp6781;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h11d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_176 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_176 <= w_sys_tmp6856;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h123: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_177 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_177 <= w_sys_tmp6931;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h129: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_178 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_178 <= w_sys_tmp7006;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp2194[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_T_datain <= w_sys_tmp2197;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp2186[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_V_datain <= w_sys_tmp2189;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp2178[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_U_datain <= w_sys_tmp2181;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3758[14:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3753[14:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3747[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3742[14:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4886[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4872[14:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4862[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4857[14:0] );

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp6548[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub09_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub09_result_datain <= w_sys_tmp3732;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_datain <= w_sys_tmp4904;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub09_result_datain <= w_sys_tmp4866;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp1979[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_T_datain <= w_sys_tmp1982;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1971[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_V_datain <= w_sys_tmp1974;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1963[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_U_datain <= w_sys_tmp1966;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3718[14:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3707[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3702[14:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3713[14:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4852[14:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4867[14:0] );

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp6473[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub08_result_datain <= w_sys_tmp3692;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub08_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub08_result_datain <= w_sys_tmp4856;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp2843[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_T_datain <= w_sys_tmp2846;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp2835[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_V_datain <= w_sys_tmp2838;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp2827[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_U_datain <= w_sys_tmp2830;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp3718[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp3713[14:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5368[14:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5353[14:0] );

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp6778[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub12_result_datain <= w_sys_tmp3720;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub12_result_datain <= w_sys_tmp5357;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp896[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_datain <= w_sys_tmp899;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp888[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_V_datain <= w_sys_tmp891;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp880[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_datain <= w_sys_tmp883;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3810[14:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3816[14:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3898[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3893[14:0] );

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp6088[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub03_result_datain <= w_sys_tmp3812;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub03_result_datain <= w_sys_tmp3902;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp681[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_datain <= w_sys_tmp684;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp673[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_V_datain <= w_sys_tmp676;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp665[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_datain <= w_sys_tmp668;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3770[14:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3776[14:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3874[14:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3903[14:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3889[14:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3879[14:0] );

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp6013[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub02_result_datain <= w_sys_tmp3772;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub02_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub02_result_datain <= w_sys_tmp3854;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp2624[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_T_datain <= w_sys_tmp2627;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp2616[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_V_datain <= w_sys_tmp2619;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp2608[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_U_datain <= w_sys_tmp2611;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3838[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3822[14:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3827[14:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3833[14:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4900[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4895[14:0] );

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp6698[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub11_result_datain <= w_sys_tmp3812;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub11_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub11_result_datain <= w_sys_tmp4904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3273[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_T_datain <= w_sys_tmp3276;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp3265[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_V_datain <= w_sys_tmp3268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp3257[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_U_datain <= w_sys_tmp3260;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp3798[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp3793[14:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5392[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5377[14:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5382[14:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp5406[14:0] );

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp6928[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub14_result_datain <= w_sys_tmp3800;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub14_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub14_result_datain <= w_sys_tmp5357;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp466[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_datain <= w_sys_tmp469;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp458[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_V_datain <= w_sys_tmp461;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp450[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_datain <= w_sys_tmp453;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3730[14:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3736[14:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3860[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3870[14:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3884[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3855[14:0] );

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp5938[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub01_result_datain <= w_sys_tmp3732;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub01_result_datain <= w_sys_tmp3902;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub01_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub01_result_datain <= w_sys_tmp3864;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3058[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_T_datain <= w_sys_tmp3061;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp3050[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_V_datain <= w_sys_tmp3053;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp3042[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_U_datain <= w_sys_tmp3045;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp3758[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp3753[14:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5387[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5358[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5373[14:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5363[14:0] );

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp6853[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub13_result_datain <= w_sys_tmp3760;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_datain <= w_sys_tmp5405;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub13_result_datain <= w_sys_tmp5367;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub13_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp251[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_datain <= w_sys_tmp254;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp243[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_V_datain <= w_sys_tmp246;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp235[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_datain <= w_sys_tmp238;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3696[14:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3690[14:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3850[14:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3865[14:0] );

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp5863[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_datain <= w_sys_tmp3692;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_datain <= w_sys_tmp3854;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp1760[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_datain <= w_sys_tmp1763;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1752[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_V_datain <= w_sys_tmp1755;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1744[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_datain <= w_sys_tmp1747;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3822[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3810[14:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3827[14:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3816[14:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4399[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4394[14:0] );

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp6393[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub07_result_datain <= w_sys_tmp3818;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub07_result_datain <= r_sys_tmp2_float;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub07_result_datain <= w_sys_tmp4403;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp1545[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_datain <= w_sys_tmp1548;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1537[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_V_datain <= w_sys_tmp1540;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1529[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_datain <= w_sys_tmp1532;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3770[14:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3787[14:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3776[14:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3782[14:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4390[14:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4380[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4375[14:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4404[14:0] );

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp6318[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub06_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub06_result_datain <= w_sys_tmp3778;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub06_result_datain <= w_sys_tmp4355;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub06_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3488[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_T_datain <= w_sys_tmp3491;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp3480[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_V_datain <= w_sys_tmp3483;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp3472[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_U_datain <= w_sys_tmp3475;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3838[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3833[14:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5401[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5396[14:0] );

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp7003[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub15_result_datain <= w_sys_tmp3840;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub15_result_datain <= w_sys_tmp5405;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp1330[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_datain <= w_sys_tmp1333;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1322[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_V_datain <= w_sys_tmp1325;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1314[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_datain <= w_sys_tmp1317;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3730[14:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3747[14:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3736[14:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3742[14:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4385[14:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4361[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4371[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4356[14:0] );

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp6243[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub05_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub05_result_datain <= w_sys_tmp3738;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub05_result_datain <= w_sys_tmp4365;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub05_result_datain <= w_sys_tmp4403;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub05_result_datain <= r_sys_tmp2_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1115[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_datain <= w_sys_tmp1118;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1107[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_V_datain <= w_sys_tmp1110;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1099[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_datain <= w_sys_tmp1102;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3707[14:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3702[14:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3696[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3690[14:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4366[14:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4351[14:0] );

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp6168[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub04_result_datain <= w_sys_tmp3698;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub04_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_datain <= w_sys_tmp4355;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp2409[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_T_datain <= w_sys_tmp2412;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp2401[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_V_datain <= w_sys_tmp2404;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp2393[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_U_datain <= w_sys_tmp2396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3798[14:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3793[14:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3787[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3782[14:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4891[14:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4905[14:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4881[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4876[14:0] );

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp6623[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub10_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub10_result_datain <= w_sys_tmp3772;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub10_result_datain <= w_sys_tmp4856;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub10_result_datain <= r_sys_tmp2_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h19)) begin
										r_sys_tmp2_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp2_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h17)) begin
										r_sys_tmp3_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp3_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h19)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp4_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
