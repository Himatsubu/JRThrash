/*
TimeStamp:	2016/11/9		15:13
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	output signed  [31:0] o_run_return	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [31:0] r_sys_run_return;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 1:0] r_sys_run_stage;
	reg         [ 3:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 1:0] w_sys_run_stage_p1;
	wire        [ 3:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_3;
	reg  signed [31:0] r_run_j_4;
	reg  signed [31:0] r_run_n_5;
	reg  signed [31:0] r_run_mx_6;
	reg  signed [31:0] r_run_my_7;
	reg  signed [31:0] r_run_nlast_8;
	reg         [31:0] r_run_dx_9;
	reg         [31:0] r_run_dy_10;
	reg         [31:0] r_run_r1_11;
	reg         [31:0] r_run_r2_12;
	reg         [31:0] r_run_dt_13;
	reg  signed [31:0] r_run_copy0_j_14;
	reg  signed [31:0] r_run_copy0_j_15;
	reg  signed [31:0] r_run_copy0_j_16;
	reg  signed [31:0] r_run_copy0_j_17;
	reg  signed [31:0] r_run_copy0_j_18;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [13:0] w_sub01_u_addr;
	reg  signed [13:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [13:0] w_sub01_result_addr;
	reg  signed [13:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [13:0] w_sub00_u_addr;
	reg  signed [13:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [13:0] w_sub00_result_addr;
	reg  signed [13:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire               w_sys_tmp8;
	wire               w_sys_tmp9;
	wire signed [31:0] w_sys_tmp10;
	wire               w_sys_tmp11;
	wire               w_sys_tmp12;
	wire signed [31:0] w_sys_tmp15;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire        [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire               w_sys_tmp56;
	wire               w_sys_tmp57;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp61;
	wire signed [31:0] w_sys_tmp62;
	wire        [31:0] w_sys_tmp63;
	wire signed [31:0] w_sys_tmp65;
	wire signed [31:0] w_sys_tmp66;
	wire        [31:0] w_sys_tmp67;
	wire signed [31:0] w_sys_tmp68;
	wire               w_sys_tmp69;
	wire               w_sys_tmp70;
	wire signed [31:0] w_sys_tmp71;
	wire signed [31:0] w_sys_tmp74;
	wire signed [31:0] w_sys_tmp75;
	wire signed [31:0] w_sys_tmp76;
	wire        [31:0] w_sys_tmp77;
	wire signed [31:0] w_sys_tmp79;
	wire signed [31:0] w_sys_tmp80;
	wire        [31:0] w_sys_tmp83;
	wire signed [31:0] w_sys_tmp84;
	wire signed [31:0] w_sys_tmp85;
	wire               w_sys_tmp164;
	wire               w_sys_tmp165;
	wire signed [31:0] w_sys_tmp166;
	wire signed [31:0] w_sys_tmp167;
	wire               w_sys_tmp168;
	wire               w_sys_tmp169;
	wire signed [31:0] w_sys_tmp170;
	wire signed [31:0] w_sys_tmp173;
	wire signed [31:0] w_sys_tmp174;
	wire signed [31:0] w_sys_tmp175;
	wire        [31:0] w_sys_tmp176;
	wire signed [31:0] w_sys_tmp177;
	wire signed [31:0] w_sys_tmp178;
	wire signed [31:0] w_sys_tmp180;
	wire signed [31:0] w_sys_tmp181;
	wire signed [31:0] w_sys_tmp242;
	wire               w_sys_tmp243;
	wire               w_sys_tmp244;
	wire signed [31:0] w_sys_tmp245;
	wire signed [31:0] w_sys_tmp248;
	wire signed [31:0] w_sys_tmp249;
	wire signed [31:0] w_sys_tmp250;
	wire signed [31:0] w_sys_tmp251;
	wire signed [31:0] w_sys_tmp252;
	wire        [31:0] w_sys_tmp253;
	wire signed [31:0] w_sys_tmp254;
	wire signed [31:0] w_sys_tmp255;
	wire signed [31:0] w_sys_tmp257;
	wire signed [31:0] w_sys_tmp258;
	wire               w_sys_tmp331;
	wire               w_sys_tmp332;
	wire signed [31:0] w_sys_tmp333;
	wire               w_sys_tmp334;
	wire               w_sys_tmp335;
	wire signed [31:0] w_sys_tmp336;
	wire signed [31:0] w_sys_tmp339;
	wire signed [31:0] w_sys_tmp340;
	wire        [31:0] w_sys_tmp341;
	wire signed [31:0] w_sys_tmp342;
	wire signed [31:0] w_sys_tmp343;
	wire signed [31:0] w_sys_tmp345;
	wire signed [31:0] w_sys_tmp346;
	wire        [31:0] w_sys_tmp347;
	wire signed [31:0] w_sys_tmp348;
	wire signed [31:0] w_sys_tmp349;
	wire signed [31:0] w_sys_tmp350;
	wire signed [31:0] w_sys_tmp351;
	wire               w_sys_tmp352;
	wire               w_sys_tmp353;
	wire signed [31:0] w_sys_tmp354;
	wire signed [31:0] w_sys_tmp355;
	wire signed [31:0] w_sys_tmp356;
	wire               w_sys_tmp357;
	wire               w_sys_tmp358;
	wire signed [31:0] w_sys_tmp359;
	wire signed [31:0] w_sys_tmp362;
	wire signed [31:0] w_sys_tmp363;
	wire signed [31:0] w_sys_tmp364;
	wire        [31:0] w_sys_tmp365;
	wire signed [31:0] w_sys_tmp366;
	wire signed [31:0] w_sys_tmp367;
	wire signed [31:0] w_sys_tmp369;
	wire signed [31:0] w_sys_tmp370;
	wire signed [31:0] w_sys_tmp431;
	wire               w_sys_tmp432;
	wire               w_sys_tmp433;
	wire signed [31:0] w_sys_tmp434;
	wire signed [31:0] w_sys_tmp437;
	wire signed [31:0] w_sys_tmp438;
	wire signed [31:0] w_sys_tmp439;
	wire        [31:0] w_sys_tmp440;
	wire signed [31:0] w_sys_tmp441;
	wire signed [31:0] w_sys_tmp442;
	wire signed [31:0] w_sys_tmp443;
	wire signed [31:0] w_sys_tmp444;
	wire signed [31:0] w_sys_tmp446;
	wire signed [31:0] w_sys_tmp447;
	wire        [31:0] w_sys_tmp520;
	wire signed [31:0] w_sys_tmp521;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign o_run_return = r_sys_run_return;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 2'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 4'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 14'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 14'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 14'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 14'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = 32'h3c000000;
	assign w_sys_tmp5 = 32'h3ba3d70a;
	assign w_sys_tmp6 = 32'h42a3d70a;
	assign w_sys_tmp8 = ( !w_sys_tmp9 );
	assign w_sys_tmp9 = (r_run_my_7 < r_run_k_3);
	assign w_sys_tmp10 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp11 = ( !w_sys_tmp12 );
	assign w_sys_tmp12 = (r_run_mx_6 < r_run_j_4);
	assign w_sys_tmp15 = (w_sys_tmp16 + r_run_k_3);
	assign w_sys_tmp16 = (r_run_j_4 * w_sys_tmp17);
	assign w_sys_tmp17 = 32'sh00000081;
	assign w_sys_tmp18 = 32'h0;
	assign w_sys_tmp19 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp56 = ( !w_sys_tmp57 );
	assign w_sys_tmp57 = (w_sys_tmp58 < r_run_k_3);
	assign w_sys_tmp58 = 32'sh00000081;
	assign w_sys_tmp61 = (w_sys_tmp62 + r_run_k_3);
	assign w_sys_tmp62 = 32'sh00000081;
	assign w_sys_tmp63 = 32'h3f000000;
	assign w_sys_tmp65 = (w_sys_tmp66 + r_run_k_3);
	assign w_sys_tmp66 = 32'sh00004101;
	assign w_sys_tmp67 = 32'h0;
	assign w_sys_tmp68 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp69 = ( !w_sys_tmp70 );
	assign w_sys_tmp70 = (w_sys_tmp71 < r_run_j_4);
	assign w_sys_tmp71 = 32'sh00000081;
	assign w_sys_tmp74 = (w_sys_tmp75 + w_sys_intOne);
	assign w_sys_tmp75 = (r_run_j_4 * w_sys_tmp76);
	assign w_sys_tmp76 = 32'sh00000081;
	assign w_sys_tmp77 = 32'h3f800000;
	assign w_sys_tmp79 = (w_sys_tmp80 + w_sys_tmp76);
	assign w_sys_tmp80 = (r_run_copy0_j_14 * w_sys_tmp76);
	assign w_sys_tmp83 = 32'h0;
	assign w_sys_tmp84 = (r_run_copy0_j_14 + w_sys_intOne);
	assign w_sys_tmp85 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp164 = ( !w_sys_tmp165 );
	assign w_sys_tmp165 = (w_sys_tmp166 < r_run_k_3);
	assign w_sys_tmp166 = 32'sh00000081;
	assign w_sys_tmp167 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp168 = ( !w_sys_tmp169 );
	assign w_sys_tmp169 = (w_sys_tmp170 < r_run_j_4);
	assign w_sys_tmp170 = 32'sh00000041;
	assign w_sys_tmp173 = (w_sys_tmp174 + r_run_k_3);
	assign w_sys_tmp174 = (r_run_j_4 * w_sys_tmp175);
	assign w_sys_tmp175 = 32'sh00000081;
	assign w_sys_tmp176 = w_fld_u_0_dataout_1;
	assign w_sys_tmp177 = (w_sys_tmp178 + r_run_k_3);
	assign w_sys_tmp178 = (r_run_copy0_j_15 * w_sys_tmp175);
	assign w_sys_tmp180 = (r_run_copy0_j_15 + w_sys_intOne);
	assign w_sys_tmp181 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp242 = 32'sh00000040;
	assign w_sys_tmp243 = ( !w_sys_tmp244 );
	assign w_sys_tmp244 = (w_sys_tmp245 < r_run_j_4);
	assign w_sys_tmp245 = 32'sh00000081;
	assign w_sys_tmp248 = (w_sys_tmp249 + r_run_k_3);
	assign w_sys_tmp249 = (w_sys_tmp250 * w_sys_tmp252);
	assign w_sys_tmp250 = (r_run_j_4 - w_sys_tmp251);
	assign w_sys_tmp251 = 32'sh0000003f;
	assign w_sys_tmp252 = 32'sh00000081;
	assign w_sys_tmp253 = w_fld_u_0_dataout_1;
	assign w_sys_tmp254 = (w_sys_tmp255 + r_run_k_3);
	assign w_sys_tmp255 = (r_run_copy0_j_16 * w_sys_tmp252);
	assign w_sys_tmp257 = (r_run_copy0_j_16 + w_sys_intOne);
	assign w_sys_tmp258 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp331 = ( !w_sys_tmp332 );
	assign w_sys_tmp332 = (r_run_nlast_8 < r_run_n_5);
	assign w_sys_tmp333 = (r_run_n_5 + w_sys_intOne);
	assign w_sys_tmp334 = ( !w_sys_tmp335 );
	assign w_sys_tmp335 = (w_sys_tmp336 < r_run_k_3);
	assign w_sys_tmp336 = 32'sh00000081;
	assign w_sys_tmp339 = (w_sys_tmp340 + r_run_k_3);
	assign w_sys_tmp340 = 32'sh00002040;
	assign w_sys_tmp341 = w_sub01_result_dataout;
	assign w_sys_tmp342 = (w_sys_tmp343 + r_run_k_3);
	assign w_sys_tmp343 = 32'sh00000081;
	assign w_sys_tmp345 = (w_sys_tmp346 + r_run_k_3);
	assign w_sys_tmp346 = 32'sh00000102;
	assign w_sys_tmp347 = w_sub00_result_dataout;
	assign w_sys_tmp348 = (w_sys_tmp349 + r_run_k_3);
	assign w_sys_tmp349 = 32'sh000020c1;
	assign w_sys_tmp350 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp351 = 32'sh00000002;
	assign w_sys_tmp352 = ( !w_sys_tmp353 );
	assign w_sys_tmp353 = (w_sys_tmp354 < r_run_k_3);
	assign w_sys_tmp354 = 32'sh00000080;
	assign w_sys_tmp355 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp356 = 32'sh00000002;
	assign w_sys_tmp357 = ( !w_sys_tmp358 );
	assign w_sys_tmp358 = (w_sys_tmp359 < r_run_j_4);
	assign w_sys_tmp359 = 32'sh00000040;
	assign w_sys_tmp362 = (w_sys_tmp363 + r_run_k_3);
	assign w_sys_tmp363 = (r_run_j_4 * w_sys_tmp364);
	assign w_sys_tmp364 = 32'sh00000081;
	assign w_sys_tmp365 = w_sub00_result_dataout;
	assign w_sys_tmp366 = (w_sys_tmp367 + r_run_k_3);
	assign w_sys_tmp367 = (r_run_copy0_j_17 * w_sys_tmp364);
	assign w_sys_tmp369 = (r_run_copy0_j_17 + w_sys_intOne);
	assign w_sys_tmp370 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp431 = 32'sh00000041;
	assign w_sys_tmp432 = ( !w_sys_tmp433 );
	assign w_sys_tmp433 = (w_sys_tmp434 < r_run_j_4);
	assign w_sys_tmp434 = 32'sh00000080;
	assign w_sys_tmp437 = (w_sys_tmp438 + r_run_k_3);
	assign w_sys_tmp438 = (r_run_j_4 * w_sys_tmp439);
	assign w_sys_tmp439 = 32'sh00000081;
	assign w_sys_tmp440 = w_sub01_result_dataout;
	assign w_sys_tmp441 = (w_sys_tmp442 + r_run_k_3);
	assign w_sys_tmp442 = (w_sys_tmp443 * w_sys_tmp439);
	assign w_sys_tmp443 = (r_run_copy0_j_18 - w_sys_tmp444);
	assign w_sys_tmp444 = 32'sh0000003f;
	assign w_sys_tmp446 = (r_run_copy0_j_18 + w_sys_intOne);
	assign w_sys_tmp447 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp520 = w_fld_u_0_dataout_1;
	assign w_sys_tmp521 = 32'sh00000104;


	subunder
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	subup
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_return <= 32'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4a: begin
							r_sys_run_return <= r_sys_tmp0_float;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h6)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp56) ? 7'h13 : 7'h15);

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp69) ? 7'h19 : 7'h1b);

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'hd)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp164) ? 7'h20 : 7'h2c);

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp168) ? 7'h24 : 7'h26);

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp243) ? 7'h2a : 7'h1d);

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp331) ? 7'h30 : 7'h3a);

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_phase <= 7'h32;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_phase <= 7'h34;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h35;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp334) ? 7'h38 : 7'h2e);

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sys_run_phase <= 7'h35;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h3b;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp352) ? 7'h3f : 7'h4b);

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h3b;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h40;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp357) ? 7'h43 : 7'h45);

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_phase <= 7'h40;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= 7'h46;

									end
								end

							endcase
						end

						7'h46: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp432) ? 7'h49 : 7'h3c);

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_phase <= 7'h46;

									end
								end

							endcase
						end

						7'h4a: begin
							r_sys_run_phase <= 7'h4d;
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sys_run_phase <= 7'h4a;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h6)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'hd)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h46: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h6)) begin
										r_sys_run_step <= 4'h0;

									end
									else
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'hd)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_step <= 4'h0;

									end
									else
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_step <= 4'h0;

									end
									else
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_step <= 4'h0;

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_step <= 4'h0;

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_step <= 4'h0;

									end
									else
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sys_run_step <= 4'h0;

									end
									else
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h1)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_step <= 4'h0;

									end
									else
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h46: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h8)) begin
										r_sys_run_step <= 4'h0;

									end
									else
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h1)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==4'h2)) begin
										r_sys_run_step <= 4'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h4d: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp15[14:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp61[14:0] );

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp65[14:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h3) || (r_sys_run_step==4'h5) || (r_sys_run_step==4'h7) || (r_sys_run_step==4'h9) || (r_sys_run_step==4'hb) || (r_sys_run_step==4'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp79[14:0] );

									end
									else
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h2) || (r_sys_run_step==4'h4) || (r_sys_run_step==4'h6) || (r_sys_run_step==4'h8) || (r_sys_run_step==4'ha) || (r_sys_run_step==4'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp74[14:0] );

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp177[14:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp254[14:0] );

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp362[14:0] );

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp437[14:0] );

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp521[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp63;

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp67;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h3) || (r_sys_run_step==4'h5) || (r_sys_run_step==4'h7) || (r_sys_run_step==4'h9) || (r_sys_run_step==4'hb) || (r_sys_run_step==4'hd)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp83;

									end
									else
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h2) || (r_sys_run_step==4'h4) || (r_sys_run_step==4'h6) || (r_sys_run_step==4'h8) || (r_sys_run_step==4'ha) || (r_sys_run_step==4'hc)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp77;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp365;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp440;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h1)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'hd)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_tmp10;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1)) begin
										r_run_k_3 <= w_sys_tmp68;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_tmp167;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_run_k_3 <= w_sys_tmp350;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_tmp351;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_k_3 <= w_sys_tmp355;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_j_4 <= w_sys_tmp19;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0) || (r_sys_run_step==4'h2) || (r_sys_run_step==4'h4) || (r_sys_run_step==4'h6) || (r_sys_run_step==4'h8) || (r_sys_run_step==4'ha) || (r_sys_run_step==4'hc)) begin
										r_run_j_4 <= w_sys_tmp85;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_run_j_4 <= w_sys_tmp181;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_tmp242;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_run_j_4 <= w_sys_tmp258;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_tmp356;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_run_j_4 <= w_sys_tmp370;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_j_4 <= w_sys_tmp431;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_run_j_4 <= w_sys_tmp447;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_n_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_n_5 <= w_sys_tmp333;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_mx_6 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_my_7 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_nlast_8 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_dx_9 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_dy_10 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_r1_11 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_r2_12 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_dt_13 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_copy0_j_14 <= r_run_j_4;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h1) || (r_sys_run_step==4'h3) || (r_sys_run_step==4'h5) || (r_sys_run_step==4'h7) || (r_sys_run_step==4'h9) || (r_sys_run_step==4'hb) || (r_sys_run_step==4'hd)) begin
										r_run_copy0_j_14 <= w_sys_tmp84;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h20: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_copy0_j_15 <= r_run_j_4;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_copy0_j_15 <= w_sys_tmp180;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_copy0_j_16 <= r_run_j_4;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_copy0_j_16 <= w_sys_tmp257;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3f: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_copy0_j_17 <= r_run_j_4;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_copy0_j_17 <= w_sys_tmp369;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_run_copy0_j_18 <= r_run_j_4;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_run_copy0_j_18 <= w_sys_tmp446;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h30: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp248[13:0] );

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp345[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_sub01_u_datain <= w_sys_tmp253;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sub01_u_datain <= w_sys_tmp347;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp342[13:0] );

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp441[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==4'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp173[13:0] );

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp339[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_sub00_u_datain <= w_sys_tmp176;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sub00_u_datain <= w_sys_tmp341;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h2<=r_sys_run_step && r_sys_run_step<=4'h8)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp348[13:0] );

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp366[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								2'h1: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((4'h0<=r_sys_run_step && r_sys_run_step<=4'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==4'h2)) begin
										r_sys_tmp0_float <= w_sys_tmp520;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
