/*
TimeStamp:	2016/6/27		14:2
*/


module c1_test02(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 2:0] r_sys_run_stage;
	reg         [ 4:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 2:0] w_sys_run_stage_p1;
	wire        [ 4:0] w_sys_run_step_p1;
	wire signed [ 8:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [ 8:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_5;
	reg  signed [31:0] r_run_j_6;
	reg  signed [31:0] r_run_n_7;
	reg  signed [31:0] r_run_mx_8;
	reg  signed [31:0] r_run_my_9;
	reg  signed [31:0] r_run_nlast_10;
	reg         [31:0] r_run_dx_11;
	reg         [31:0] r_run_dy_12;
	reg  signed [31:0] r_run_copy0_j_13;
	reg  signed [31:0] r_run_copy1_j_14;
	reg  signed [31:0] r_run_copy2_j_15;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 8:0] w_sub03_u_addr;
	reg  signed [ 8:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [ 8:0] w_sub03_result_addr;
	reg  signed [ 8:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 8:0] w_sub02_u_addr;
	reg  signed [ 8:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [ 8:0] w_sub02_result_addr;
	reg  signed [ 8:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 9:0] w_sub01_u_addr;
	reg  signed [ 9:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [ 9:0] w_sub01_result_addr;
	reg  signed [ 9:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 8:0] w_sub00_u_addr;
	reg  signed [ 8:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [ 8:0] w_sub00_result_addr;
	reg  signed [ 8:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire               w_sys_tmp5;
	wire               w_sys_tmp6;
	wire signed [31:0] w_sys_tmp7;
	wire               w_sys_tmp8;
	wire               w_sys_tmp9;
	wire signed [31:0] w_sys_tmp12;
	wire signed [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire        [31:0] w_sys_tmp15;
	wire signed [31:0] w_sys_tmp16;
	wire               w_sys_tmp53;
	wire               w_sys_tmp54;
	wire signed [31:0] w_sys_tmp55;
	wire               w_sys_tmp56;
	wire               w_sys_tmp57;
	wire signed [31:0] w_sys_tmp60;
	wire signed [31:0] w_sys_tmp61;
	wire        [31:0] w_sys_tmp62;
	wire signed [31:0] w_sys_tmp64;
	wire signed [31:0] w_sys_tmp65;
	wire        [31:0] w_sys_tmp67;
	wire signed [31:0] w_sys_tmp69;
	wire signed [31:0] w_sys_tmp70;
	wire        [31:0] w_sys_tmp72;
	wire signed [31:0] w_sys_tmp74;
	wire signed [31:0] w_sys_tmp75;
	wire signed [31:0] w_sys_tmp78;
	wire signed [31:0] w_sys_tmp79;
	wire signed [31:0] w_sys_tmp80;
	wire signed [31:0] w_sys_tmp81;
	wire signed [31:0] w_sys_tmp220;
	wire               w_sys_tmp221;
	wire               w_sys_tmp222;
	wire signed [31:0] w_sys_tmp225;
	wire signed [31:0] w_sys_tmp226;
	wire        [31:0] w_sys_tmp227;
	wire signed [31:0] w_sys_tmp231;
	wire signed [31:0] w_sys_tmp232;
	wire signed [31:0] w_sys_tmp237;
	wire signed [31:0] w_sys_tmp238;
	wire signed [31:0] w_sys_tmp243;
	wire signed [31:0] w_sys_tmp244;
	wire signed [31:0] w_sys_tmp249;
	wire signed [31:0] w_sys_tmp250;
	wire signed [31:0] w_sys_tmp255;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp261;
	wire signed [31:0] w_sys_tmp262;
	wire signed [31:0] w_sys_tmp267;
	wire signed [31:0] w_sys_tmp268;
	wire signed [31:0] w_sys_tmp273;
	wire signed [31:0] w_sys_tmp274;
	wire signed [31:0] w_sys_tmp279;
	wire signed [31:0] w_sys_tmp280;
	wire signed [31:0] w_sys_tmp285;
	wire signed [31:0] w_sys_tmp286;
	wire signed [31:0] w_sys_tmp291;
	wire signed [31:0] w_sys_tmp292;
	wire signed [31:0] w_sys_tmp297;
	wire signed [31:0] w_sys_tmp298;
	wire signed [31:0] w_sys_tmp303;
	wire signed [31:0] w_sys_tmp304;
	wire signed [31:0] w_sys_tmp309;
	wire signed [31:0] w_sys_tmp310;
	wire signed [31:0] w_sys_tmp315;
	wire signed [31:0] w_sys_tmp316;
	wire signed [31:0] w_sys_tmp321;
	wire signed [31:0] w_sys_tmp322;
	wire signed [31:0] w_sys_tmp327;
	wire signed [31:0] w_sys_tmp328;
	wire signed [31:0] w_sys_tmp333;
	wire signed [31:0] w_sys_tmp334;
	wire signed [31:0] w_sys_tmp339;
	wire signed [31:0] w_sys_tmp340;
	wire signed [31:0] w_sys_tmp345;
	wire signed [31:0] w_sys_tmp346;
	wire signed [31:0] w_sys_tmp362;
	wire               w_sys_tmp363;
	wire               w_sys_tmp364;
	wire signed [31:0] w_sys_tmp365;
	wire signed [31:0] w_sys_tmp368;
	wire signed [31:0] w_sys_tmp369;
	wire        [31:0] w_sys_tmp370;
	wire signed [31:0] w_sys_tmp374;
	wire signed [31:0] w_sys_tmp375;
	wire signed [31:0] w_sys_tmp380;
	wire signed [31:0] w_sys_tmp381;
	wire signed [31:0] w_sys_tmp386;
	wire signed [31:0] w_sys_tmp387;
	wire signed [31:0] w_sys_tmp392;
	wire signed [31:0] w_sys_tmp393;
	wire signed [31:0] w_sys_tmp398;
	wire signed [31:0] w_sys_tmp399;
	wire signed [31:0] w_sys_tmp404;
	wire signed [31:0] w_sys_tmp405;
	wire signed [31:0] w_sys_tmp410;
	wire signed [31:0] w_sys_tmp411;
	wire signed [31:0] w_sys_tmp416;
	wire signed [31:0] w_sys_tmp417;
	wire signed [31:0] w_sys_tmp422;
	wire signed [31:0] w_sys_tmp423;
	wire signed [31:0] w_sys_tmp428;
	wire signed [31:0] w_sys_tmp429;
	wire signed [31:0] w_sys_tmp434;
	wire signed [31:0] w_sys_tmp435;
	wire signed [31:0] w_sys_tmp440;
	wire signed [31:0] w_sys_tmp441;
	wire signed [31:0] w_sys_tmp446;
	wire signed [31:0] w_sys_tmp447;
	wire signed [31:0] w_sys_tmp452;
	wire signed [31:0] w_sys_tmp453;
	wire signed [31:0] w_sys_tmp458;
	wire signed [31:0] w_sys_tmp459;
	wire signed [31:0] w_sys_tmp464;
	wire signed [31:0] w_sys_tmp465;
	wire signed [31:0] w_sys_tmp470;
	wire signed [31:0] w_sys_tmp471;
	wire signed [31:0] w_sys_tmp476;
	wire signed [31:0] w_sys_tmp477;
	wire signed [31:0] w_sys_tmp482;
	wire signed [31:0] w_sys_tmp483;
	wire signed [31:0] w_sys_tmp488;
	wire signed [31:0] w_sys_tmp489;
	wire signed [31:0] w_sys_tmp505;
	wire signed [31:0] w_sys_tmp506;
	wire               w_sys_tmp507;
	wire               w_sys_tmp508;
	wire signed [31:0] w_sys_tmp509;
	wire signed [31:0] w_sys_tmp512;
	wire signed [31:0] w_sys_tmp513;
	wire        [31:0] w_sys_tmp514;
	wire signed [31:0] w_sys_tmp515;
	wire signed [31:0] w_sys_tmp516;
	wire signed [31:0] w_sys_tmp517;
	wire signed [31:0] w_sys_tmp519;
	wire signed [31:0] w_sys_tmp520;
	wire signed [31:0] w_sys_tmp526;
	wire signed [31:0] w_sys_tmp527;
	wire signed [31:0] w_sys_tmp533;
	wire signed [31:0] w_sys_tmp534;
	wire signed [31:0] w_sys_tmp540;
	wire signed [31:0] w_sys_tmp541;
	wire signed [31:0] w_sys_tmp547;
	wire signed [31:0] w_sys_tmp548;
	wire signed [31:0] w_sys_tmp554;
	wire signed [31:0] w_sys_tmp555;
	wire signed [31:0] w_sys_tmp561;
	wire signed [31:0] w_sys_tmp562;
	wire signed [31:0] w_sys_tmp568;
	wire signed [31:0] w_sys_tmp569;
	wire signed [31:0] w_sys_tmp575;
	wire signed [31:0] w_sys_tmp576;
	wire signed [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp581;
	wire signed [31:0] w_sys_tmp585;
	wire signed [31:0] w_sys_tmp586;
	wire signed [31:0] w_sys_tmp590;
	wire signed [31:0] w_sys_tmp591;
	wire signed [31:0] w_sys_tmp595;
	wire signed [31:0] w_sys_tmp596;
	wire signed [31:0] w_sys_tmp600;
	wire signed [31:0] w_sys_tmp601;
	wire signed [31:0] w_sys_tmp605;
	wire signed [31:0] w_sys_tmp606;
	wire signed [31:0] w_sys_tmp610;
	wire signed [31:0] w_sys_tmp611;
	wire signed [31:0] w_sys_tmp615;
	wire signed [31:0] w_sys_tmp616;
	wire signed [31:0] w_sys_tmp620;
	wire signed [31:0] w_sys_tmp621;
	wire signed [31:0] w_sys_tmp624;
	wire signed [31:0] w_sys_tmp625;
	wire               w_sys_tmp626;
	wire               w_sys_tmp627;
	wire signed [31:0] w_sys_tmp628;
	wire signed [31:0] w_sys_tmp631;
	wire signed [31:0] w_sys_tmp632;
	wire        [31:0] w_sys_tmp633;
	wire signed [31:0] w_sys_tmp637;
	wire signed [31:0] w_sys_tmp638;
	wire signed [31:0] w_sys_tmp643;
	wire signed [31:0] w_sys_tmp644;
	wire signed [31:0] w_sys_tmp649;
	wire signed [31:0] w_sys_tmp650;
	wire signed [31:0] w_sys_tmp655;
	wire signed [31:0] w_sys_tmp656;
	wire signed [31:0] w_sys_tmp661;
	wire signed [31:0] w_sys_tmp662;
	wire signed [31:0] w_sys_tmp667;
	wire signed [31:0] w_sys_tmp668;
	wire signed [31:0] w_sys_tmp673;
	wire signed [31:0] w_sys_tmp674;
	wire signed [31:0] w_sys_tmp679;
	wire signed [31:0] w_sys_tmp680;
	wire signed [31:0] w_sys_tmp685;
	wire signed [31:0] w_sys_tmp686;
	wire signed [31:0] w_sys_tmp690;
	wire signed [31:0] w_sys_tmp691;
	wire signed [31:0] w_sys_tmp695;
	wire signed [31:0] w_sys_tmp696;
	wire signed [31:0] w_sys_tmp700;
	wire signed [31:0] w_sys_tmp701;
	wire signed [31:0] w_sys_tmp705;
	wire signed [31:0] w_sys_tmp706;
	wire signed [31:0] w_sys_tmp710;
	wire signed [31:0] w_sys_tmp711;
	wire signed [31:0] w_sys_tmp715;
	wire signed [31:0] w_sys_tmp716;
	wire signed [31:0] w_sys_tmp720;
	wire signed [31:0] w_sys_tmp721;
	wire signed [31:0] w_sys_tmp725;
	wire signed [31:0] w_sys_tmp726;
	wire signed [31:0] w_sys_tmp730;
	wire signed [31:0] w_sys_tmp731;
	wire signed [31:0] w_sys_tmp734;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 3'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 5'h1);
	assign w_fld_u_0_addr_0 = 9'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 9'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 9'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 9'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 9'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 10'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 10'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 9'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 9'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000015;
	assign w_sys_tmp3 = 32'h3d4ccccd;
	assign w_sys_tmp5 = ( !w_sys_tmp6 );
	assign w_sys_tmp6 = (r_run_my_9 < r_run_k_5);
	assign w_sys_tmp7 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp8 = ( !w_sys_tmp9 );
	assign w_sys_tmp9 = (r_run_mx_8 < r_run_j_6);
	assign w_sys_tmp12 = (w_sys_tmp13 + r_run_k_5);
	assign w_sys_tmp13 = (r_run_j_6 * w_sys_tmp14);
	assign w_sys_tmp14 = 32'sh00000015;
	assign w_sys_tmp15 = 32'h0;
	assign w_sys_tmp16 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp53 = ( !w_sys_tmp54 );
	assign w_sys_tmp54 = (r_run_nlast_10 < r_run_n_7);
	assign w_sys_tmp55 = (r_run_n_7 + w_sys_intOne);
	assign w_sys_tmp56 = ( !w_sys_tmp57 );
	assign w_sys_tmp57 = (r_run_my_9 < r_run_j_6);
	assign w_sys_tmp60 = (w_sys_tmp61 + r_run_j_6);
	assign w_sys_tmp61 = 32'sh00000015;
	assign w_sys_tmp62 = 32'h3f000000;
	assign w_sys_tmp64 = (w_sys_tmp65 + r_run_copy2_j_15);
	assign w_sys_tmp65 = (r_run_mx_8 * w_sys_tmp61);
	assign w_sys_tmp67 = 32'h0;
	assign w_sys_tmp69 = (w_sys_tmp70 + w_sys_intOne);
	assign w_sys_tmp70 = (r_run_copy1_j_14 * w_sys_tmp61);
	assign w_sys_tmp72 = 32'h3f800000;
	assign w_sys_tmp74 = (w_sys_tmp75 + r_run_my_9);
	assign w_sys_tmp75 = (r_run_copy0_j_13 * w_sys_tmp61);
	assign w_sys_tmp78 = (r_run_copy0_j_13 + w_sys_intOne);
	assign w_sys_tmp79 = (r_run_copy1_j_14 + w_sys_intOne);
	assign w_sys_tmp80 = (r_run_copy2_j_15 + w_sys_intOne);
	assign w_sys_tmp81 = (r_run_j_6 + w_sys_intOne);
	assign w_sys_tmp220 = 32'sh0000000a;
	assign w_sys_tmp221 = ( !w_sys_tmp222 );
	assign w_sys_tmp222 = (r_run_my_9 < r_run_k_5);
	assign w_sys_tmp225 = (w_sys_tmp226 + r_run_k_5);
	assign w_sys_tmp226 = 32'sh000000d2;
	assign w_sys_tmp227 = w_fld_u_0_dataout_1;
	assign w_sys_tmp231 = (w_sys_tmp232 + r_run_k_5);
	assign w_sys_tmp232 = 32'sh000000e7;
	assign w_sys_tmp237 = (w_sys_tmp238 + r_run_k_5);
	assign w_sys_tmp238 = 32'sh000000fc;
	assign w_sys_tmp243 = (w_sys_tmp244 + r_run_k_5);
	assign w_sys_tmp244 = 32'sh00000111;
	assign w_sys_tmp249 = (w_sys_tmp250 + r_run_k_5);
	assign w_sys_tmp250 = 32'sh00000126;
	assign w_sys_tmp255 = (w_sys_tmp256 + r_run_k_5);
	assign w_sys_tmp256 = 32'sh0000013b;
	assign w_sys_tmp261 = (w_sys_tmp262 + r_run_k_5);
	assign w_sys_tmp262 = 32'sh00000150;
	assign w_sys_tmp267 = (w_sys_tmp268 + r_run_k_5);
	assign w_sys_tmp268 = 32'sh00000165;
	assign w_sys_tmp273 = (w_sys_tmp274 + r_run_k_5);
	assign w_sys_tmp274 = 32'sh0000017a;
	assign w_sys_tmp279 = (w_sys_tmp280 + r_run_k_5);
	assign w_sys_tmp280 = 32'sh0000018f;
	assign w_sys_tmp285 = (w_sys_tmp286 + r_run_k_5);
	assign w_sys_tmp286 = 32'sh000001a4;
	assign w_sys_tmp291 = (w_sys_tmp292 + r_run_k_5);
	assign w_sys_tmp292 = 32'sh000001b9;
	assign w_sys_tmp297 = (w_sys_tmp298 + r_run_k_5);
	assign w_sys_tmp298 = 32'sh00000015;
	assign w_sys_tmp303 = (w_sys_tmp304 + r_run_k_5);
	assign w_sys_tmp304 = 32'sh0000002a;
	assign w_sys_tmp309 = (w_sys_tmp310 + r_run_k_5);
	assign w_sys_tmp310 = 32'sh0000003f;
	assign w_sys_tmp315 = (w_sys_tmp316 + r_run_k_5);
	assign w_sys_tmp316 = 32'sh00000054;
	assign w_sys_tmp321 = (w_sys_tmp322 + r_run_k_5);
	assign w_sys_tmp322 = 32'sh00000069;
	assign w_sys_tmp327 = (w_sys_tmp328 + r_run_k_5);
	assign w_sys_tmp328 = 32'sh0000007e;
	assign w_sys_tmp333 = (w_sys_tmp334 + r_run_k_5);
	assign w_sys_tmp334 = 32'sh00000093;
	assign w_sys_tmp339 = (w_sys_tmp340 + r_run_k_5);
	assign w_sys_tmp340 = 32'sh000000a8;
	assign w_sys_tmp345 = (w_sys_tmp346 + r_run_k_5);
	assign w_sys_tmp346 = 32'sh000000bd;
	assign w_sys_tmp362 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp363 = ( !w_sys_tmp364 );
	assign w_sys_tmp364 = (w_sys_tmp365 < r_run_k_5);
	assign w_sys_tmp365 = 32'sh0000000b;
	assign w_sys_tmp368 = (w_sys_tmp369 + r_run_k_5);
	assign w_sys_tmp369 = 32'sh000000d2;
	assign w_sys_tmp370 = w_fld_u_0_dataout_1;
	assign w_sys_tmp374 = (w_sys_tmp375 + r_run_k_5);
	assign w_sys_tmp375 = 32'sh000000e7;
	assign w_sys_tmp380 = (w_sys_tmp381 + r_run_k_5);
	assign w_sys_tmp381 = 32'sh000000fc;
	assign w_sys_tmp386 = (w_sys_tmp387 + r_run_k_5);
	assign w_sys_tmp387 = 32'sh00000111;
	assign w_sys_tmp392 = (w_sys_tmp393 + r_run_k_5);
	assign w_sys_tmp393 = 32'sh00000126;
	assign w_sys_tmp398 = (w_sys_tmp399 + r_run_k_5);
	assign w_sys_tmp399 = 32'sh0000013b;
	assign w_sys_tmp404 = (w_sys_tmp405 + r_run_k_5);
	assign w_sys_tmp405 = 32'sh00000150;
	assign w_sys_tmp410 = (w_sys_tmp411 + r_run_k_5);
	assign w_sys_tmp411 = 32'sh00000165;
	assign w_sys_tmp416 = (w_sys_tmp417 + r_run_k_5);
	assign w_sys_tmp417 = 32'sh0000017a;
	assign w_sys_tmp422 = (w_sys_tmp423 + r_run_k_5);
	assign w_sys_tmp423 = 32'sh0000018f;
	assign w_sys_tmp428 = (w_sys_tmp429 + r_run_k_5);
	assign w_sys_tmp429 = 32'sh000001a4;
	assign w_sys_tmp434 = (w_sys_tmp435 + r_run_k_5);
	assign w_sys_tmp435 = 32'sh000001b9;
	assign w_sys_tmp440 = (w_sys_tmp441 + r_run_k_5);
	assign w_sys_tmp441 = 32'sh00000015;
	assign w_sys_tmp446 = (w_sys_tmp447 + r_run_k_5);
	assign w_sys_tmp447 = 32'sh0000002a;
	assign w_sys_tmp452 = (w_sys_tmp453 + r_run_k_5);
	assign w_sys_tmp453 = 32'sh0000003f;
	assign w_sys_tmp458 = (w_sys_tmp459 + r_run_k_5);
	assign w_sys_tmp459 = 32'sh00000054;
	assign w_sys_tmp464 = (w_sys_tmp465 + r_run_k_5);
	assign w_sys_tmp465 = 32'sh00000069;
	assign w_sys_tmp470 = (w_sys_tmp471 + r_run_k_5);
	assign w_sys_tmp471 = 32'sh0000007e;
	assign w_sys_tmp476 = (w_sys_tmp477 + r_run_k_5);
	assign w_sys_tmp477 = 32'sh00000093;
	assign w_sys_tmp482 = (w_sys_tmp483 + r_run_k_5);
	assign w_sys_tmp483 = 32'sh000000a8;
	assign w_sys_tmp488 = (w_sys_tmp489 + r_run_k_5);
	assign w_sys_tmp489 = 32'sh000000bd;
	assign w_sys_tmp505 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp506 = 32'sh00000002;
	assign w_sys_tmp507 = ( !w_sys_tmp508 );
	assign w_sys_tmp508 = (w_sys_tmp509 < r_run_k_5);
	assign w_sys_tmp509 = 32'sh0000000a;
	assign w_sys_tmp512 = (w_sys_tmp513 + r_run_k_5);
	assign w_sys_tmp513 = 32'sh0000002a;
	assign w_sys_tmp514 = w_sub00_result_dataout;
	assign w_sys_tmp515 = (w_sys_tmp516 + r_run_k_5);
	assign w_sys_tmp516 = (r_run_j_6 * w_sys_tmp517);
	assign w_sys_tmp517 = 32'sh00000015;
	assign w_sys_tmp519 = (w_sys_tmp520 + r_run_k_5);
	assign w_sys_tmp520 = 32'sh0000003f;
	assign w_sys_tmp526 = (w_sys_tmp527 + r_run_k_5);
	assign w_sys_tmp527 = 32'sh00000054;
	assign w_sys_tmp533 = (w_sys_tmp534 + r_run_k_5);
	assign w_sys_tmp534 = 32'sh00000069;
	assign w_sys_tmp540 = (w_sys_tmp541 + r_run_k_5);
	assign w_sys_tmp541 = 32'sh0000007e;
	assign w_sys_tmp547 = (w_sys_tmp548 + r_run_k_5);
	assign w_sys_tmp548 = 32'sh00000093;
	assign w_sys_tmp554 = (w_sys_tmp555 + r_run_k_5);
	assign w_sys_tmp555 = 32'sh000000a8;
	assign w_sys_tmp561 = (w_sys_tmp562 + r_run_k_5);
	assign w_sys_tmp562 = 32'sh000000bd;
	assign w_sys_tmp568 = (w_sys_tmp569 + r_run_k_5);
	assign w_sys_tmp569 = 32'sh000000d2;
	assign w_sys_tmp575 = (w_sys_tmp576 + r_run_k_5);
	assign w_sys_tmp576 = 32'sh000000e7;
	assign w_sys_tmp580 = (w_sys_tmp581 + r_run_k_5);
	assign w_sys_tmp581 = 32'sh000000fc;
	assign w_sys_tmp585 = (w_sys_tmp586 + r_run_k_5);
	assign w_sys_tmp586 = 32'sh00000111;
	assign w_sys_tmp590 = (w_sys_tmp591 + r_run_k_5);
	assign w_sys_tmp591 = 32'sh00000126;
	assign w_sys_tmp595 = (w_sys_tmp596 + r_run_k_5);
	assign w_sys_tmp596 = 32'sh0000013b;
	assign w_sys_tmp600 = (w_sys_tmp601 + r_run_k_5);
	assign w_sys_tmp601 = 32'sh00000150;
	assign w_sys_tmp605 = (w_sys_tmp606 + r_run_k_5);
	assign w_sys_tmp606 = 32'sh00000165;
	assign w_sys_tmp610 = (w_sys_tmp611 + r_run_k_5);
	assign w_sys_tmp611 = 32'sh0000017a;
	assign w_sys_tmp615 = (w_sys_tmp616 + r_run_k_5);
	assign w_sys_tmp616 = 32'sh0000018f;
	assign w_sys_tmp620 = (w_sys_tmp621 + r_run_k_5);
	assign w_sys_tmp621 = 32'sh000001a4;
	assign w_sys_tmp624 = (r_run_k_5 + w_sys_intOne);
	assign w_sys_tmp625 = 32'sh0000000b;
	assign w_sys_tmp626 = ( !w_sys_tmp627 );
	assign w_sys_tmp627 = (w_sys_tmp628 < r_run_k_5);
	assign w_sys_tmp628 = 32'sh00000014;
	assign w_sys_tmp631 = (w_sys_tmp632 + r_run_k_5);
	assign w_sys_tmp632 = 32'sh0000002a;
	assign w_sys_tmp633 = w_sub02_result_dataout;
	assign w_sys_tmp637 = (w_sys_tmp638 + r_run_k_5);
	assign w_sys_tmp638 = 32'sh0000003f;
	assign w_sys_tmp643 = (w_sys_tmp644 + r_run_k_5);
	assign w_sys_tmp644 = 32'sh00000054;
	assign w_sys_tmp649 = (w_sys_tmp650 + r_run_k_5);
	assign w_sys_tmp650 = 32'sh00000069;
	assign w_sys_tmp655 = (w_sys_tmp656 + r_run_k_5);
	assign w_sys_tmp656 = 32'sh0000007e;
	assign w_sys_tmp661 = (w_sys_tmp662 + r_run_k_5);
	assign w_sys_tmp662 = 32'sh00000093;
	assign w_sys_tmp667 = (w_sys_tmp668 + r_run_k_5);
	assign w_sys_tmp668 = 32'sh000000a8;
	assign w_sys_tmp673 = (w_sys_tmp674 + r_run_k_5);
	assign w_sys_tmp674 = 32'sh000000bd;
	assign w_sys_tmp679 = (w_sys_tmp680 + r_run_k_5);
	assign w_sys_tmp680 = 32'sh000000d2;
	assign w_sys_tmp685 = (w_sys_tmp686 + r_run_k_5);
	assign w_sys_tmp686 = 32'sh000000e7;
	assign w_sys_tmp690 = (w_sys_tmp691 + r_run_k_5);
	assign w_sys_tmp691 = 32'sh000000fc;
	assign w_sys_tmp695 = (w_sys_tmp696 + r_run_k_5);
	assign w_sys_tmp696 = 32'sh00000111;
	assign w_sys_tmp700 = (w_sys_tmp701 + r_run_k_5);
	assign w_sys_tmp701 = 32'sh00000126;
	assign w_sys_tmp705 = (w_sys_tmp706 + r_run_k_5);
	assign w_sys_tmp706 = 32'sh0000013b;
	assign w_sys_tmp710 = (w_sys_tmp711 + r_run_k_5);
	assign w_sys_tmp711 = 32'sh00000150;
	assign w_sys_tmp715 = (w_sys_tmp716 + r_run_k_5);
	assign w_sys_tmp716 = 32'sh00000165;
	assign w_sys_tmp720 = (w_sys_tmp721 + r_run_k_5);
	assign w_sys_tmp721 = 32'sh0000017a;
	assign w_sys_tmp725 = (w_sys_tmp726 + r_run_k_5);
	assign w_sys_tmp726 = 32'sh0000018f;
	assign w_sys_tmp730 = (w_sys_tmp731 + r_run_k_5);
	assign w_sys_tmp731 = 32'sh000001a4;
	assign w_sys_tmp734 = (r_run_k_5 + w_sys_intOne);


	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h35: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp53) ? 6'h14 : 6'h35);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp56) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp221) ? 6'h1e : 6'h20);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h18)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp363) ? 6'h24 : 6'h25);

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h18)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 6'h27;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_phase <= 6'h29;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp507) ? 6'h2d : 6'h2f);

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h14)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp626) ? 6'h33 : 6'h11);

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h14)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h35: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 3'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h18)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h18)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h14)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h14)) begin
										r_sys_run_stage <= 3'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==5'h1b)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h18)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h17)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h18)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h17)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h1)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h14)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h13)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sys_run_step <= 5'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h14)) begin
										r_sys_run_step <= 5'h0;

									end
									else
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h13)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h35: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp12[8:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp64[8:0] );

									end
									else
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp60[8:0] );

									end
									else
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp69[8:0] );

									end
									else
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp74[8:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp273[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp249[8:0] );

									end
									else
									if((r_sys_run_step==5'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp321[8:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp279[8:0] );

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp231[8:0] );

									end
									else
									if((r_sys_run_step==5'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp285[8:0] );

									end
									else
									if((r_sys_run_step==5'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp297[8:0] );

									end
									else
									if((r_sys_run_step==5'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp345[8:0] );

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp261[8:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp291[8:0] );

									end
									else
									if((r_sys_run_step==5'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp339[8:0] );

									end
									else
									if((r_sys_run_step==5'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp303[8:0] );

									end
									else
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp225[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp267[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp237[8:0] );

									end
									else
									if((r_sys_run_step==5'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp309[8:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp255[8:0] );

									end
									else
									if((r_sys_run_step==5'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp333[8:0] );

									end
									else
									if((r_sys_run_step==5'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp327[8:0] );

									end
									else
									if((r_sys_run_step==5'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp315[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp243[8:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp470[8:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp422[8:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp434[8:0] );

									end
									else
									if((r_sys_run_step==5'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp428[8:0] );

									end
									else
									if((r_sys_run_step==5'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp452[8:0] );

									end
									else
									if((r_sys_run_step==5'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp464[8:0] );

									end
									else
									if((r_sys_run_step==5'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp458[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp380[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp410[8:0] );

									end
									else
									if((r_sys_run_step==5'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp446[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp392[8:0] );

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp374[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp386[8:0] );

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp404[8:0] );

									end
									else
									if((r_sys_run_step==5'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp440[8:0] );

									end
									else
									if((r_sys_run_step==5'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp482[8:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp398[8:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp416[8:0] );

									end
									else
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp368[8:0] );

									end
									else
									if((r_sys_run_step==5'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp488[8:0] );

									end
									else
									if((r_sys_run_step==5'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp476[8:0] );

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==5'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp595[8:0] );

									end
									else
									if((r_sys_run_step==5'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp615[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp526[8:0] );

									end
									else
									if((r_sys_run_step==5'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp600[8:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp561[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp519[8:0] );

									end
									else
									if((r_sys_run_step==5'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp590[8:0] );

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp540[8:0] );

									end
									else
									if((r_sys_run_step==5'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp585[8:0] );

									end
									else
									if((r_sys_run_step==5'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp568[8:0] );

									end
									else
									if((r_sys_run_step==5'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp610[8:0] );

									end
									else
									if((r_sys_run_step==5'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp620[8:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp533[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp547[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp512[8:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp575[8:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp554[8:0] );

									end
									else
									if((r_sys_run_step==5'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp605[8:0] );

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp637[8:0] );

									end
									else
									if((r_sys_run_step==5'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp679[8:0] );

									end
									else
									if((r_sys_run_step==5'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp695[8:0] );

									end
									else
									if((r_sys_run_step==5'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp730[8:0] );

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp655[8:0] );

									end
									else
									if((r_sys_run_step==5'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp715[8:0] );

									end
									else
									if((r_sys_run_step==5'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp720[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp661[8:0] );

									end
									else
									if((r_sys_run_step==5'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp725[8:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp685[8:0] );

									end
									else
									if((r_sys_run_step==5'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp705[8:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp649[8:0] );

									end
									else
									if((r_sys_run_step==5'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp700[8:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp667[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp643[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp631[8:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp673[8:0] );

									end
									else
									if((r_sys_run_step==5'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp690[8:0] );

									end
									else
									if((r_sys_run_step==5'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp710[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp15;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp62;

									end
									else
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp72;

									end
									else
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h3) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h19) || (r_sys_run_step==5'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp67;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==5'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'ha)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp514;

									end
									else
									if((r_sys_run_step==5'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==5'hb) || (r_sys_run_step==5'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==5'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==5'hc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==5'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==5'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==5'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==5'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==5'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==5'hb) || (r_sys_run_step==5'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==5'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'ha)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp633;

									end
									else
									if((r_sys_run_step==5'hc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==5'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==5'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==5'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h16)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h16)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h14)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'h14)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h35: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp7;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp220;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h18)) begin
										r_run_k_5 <= w_sys_tmp362;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h18)) begin
										r_run_k_5 <= w_sys_tmp505;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp506;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h14)) begin
										r_run_k_5 <= w_sys_tmp624;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_k_5 <= w_sys_tmp625;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h14)) begin
										r_run_k_5 <= w_sys_tmp734;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h6)) begin
										r_run_j_6 <= w_sys_tmp16;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_j_6 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0) || (r_sys_run_step==5'h4) || (r_sys_run_step==5'h8) || (r_sys_run_step==5'hc) || (r_sys_run_step==5'h10) || (r_sys_run_step==5'h14) || (r_sys_run_step==5'h18)) begin
										r_run_j_6 <= w_sys_tmp81;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_n_7 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_n_7 <= w_sys_tmp55;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_mx_8 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_my_9 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_nlast_10 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_dx_11 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_dy_12 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy0_j_13 <= r_run_j_6;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3) || (r_sys_run_step==5'h7) || (r_sys_run_step==5'hb) || (r_sys_run_step==5'hf) || (r_sys_run_step==5'h13) || (r_sys_run_step==5'h17) || (r_sys_run_step==5'h1b)) begin
										r_run_copy0_j_13 <= w_sys_tmp78;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy1_j_14 <= r_run_j_6;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'h6) || (r_sys_run_step==5'ha) || (r_sys_run_step==5'he) || (r_sys_run_step==5'h12) || (r_sys_run_step==5'h16) || (r_sys_run_step==5'h1a)) begin
										r_run_copy1_j_14 <= w_sys_tmp79;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_run_copy2_j_15 <= r_run_j_6;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1) || (r_sys_run_step==5'h5) || (r_sys_run_step==5'h9) || (r_sys_run_step==5'hd) || (r_sys_run_step==5'h11) || (r_sys_run_step==5'h15) || (r_sys_run_step==5'h19)) begin
										r_run_copy2_j_15 <= w_sys_tmp80;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'ha)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp273[8:0] );

									end
									else
									if((r_sys_run_step==5'hd)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp291[8:0] );

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp249[8:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp279[8:0] );

									end
									else
									if((r_sys_run_step==5'hc)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp285[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp231[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp225[8:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp267[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp237[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp255[8:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp261[8:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp243[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'hd)) begin
										r_sub03_u_datain <= w_sys_tmp227;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'hd)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp715[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp720[8:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp725[8:0] );

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp685[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp705[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp695[8:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp730[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp700[8:0] );

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp690[8:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp710[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h9)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h15)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp339[8:0] );

									end
									else
									if((r_sys_run_step==5'h12)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp321[8:0] );

									end
									else
									if((r_sys_run_step==5'h18)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp231[8:0] );

									end
									else
									if((r_sys_run_step==5'hf)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp303[8:0] );

									end
									else
									if((r_sys_run_step==5'he)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp297[8:0] );

									end
									else
									if((r_sys_run_step==5'h17)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp225[8:0] );

									end
									else
									if((r_sys_run_step==5'h16)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp345[8:0] );

									end
									else
									if((r_sys_run_step==5'h10)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp309[8:0] );

									end
									else
									if((r_sys_run_step==5'h14)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp333[8:0] );

									end
									else
									if((r_sys_run_step==5'h13)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp327[8:0] );

									end
									else
									if((r_sys_run_step==5'h11)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp315[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'he<=r_sys_run_step && r_sys_run_step<=5'h18)) begin
										r_sub02_u_datain <= w_sys_tmp227;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'he<=r_sys_run_step && r_sys_run_step<=5'h18)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp637[8:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp679[8:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp661[8:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp649[8:0] );

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp667[8:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp643[8:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp673[8:0] );

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp631[8:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp655[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp374[9:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp404[9:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp386[9:0] );

									end
									else
									if((r_sys_run_step==5'hd)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp434[9:0] );

									end
									else
									if((r_sys_run_step==5'hb)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp422[9:0] );

									end
									else
									if((r_sys_run_step==5'hc)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp428[9:0] );

									end
									else
									if((r_sys_run_step==5'ha)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp416[9:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp398[9:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp368[9:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp410[9:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp380[9:0] );

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp392[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'hd)) begin
										r_sub01_u_datain <= w_sys_tmp370;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h2<=r_sys_run_step && r_sys_run_step<=5'hd)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp580[9:0] );

									end
									else
									if((r_sys_run_step==5'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp595[9:0] );

									end
									else
									if((r_sys_run_step==5'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp610[9:0] );

									end
									else
									if((r_sys_run_step==5'h9)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp620[9:0] );

									end
									else
									if((r_sys_run_step==5'h8)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp615[9:0] );

									end
									else
									if((r_sys_run_step==5'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp600[9:0] );

									end
									else
									if((r_sys_run_step==5'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp590[9:0] );

									end
									else
									if((r_sys_run_step==5'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp585[9:0] );

									end
									else
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp575[9:0] );

									end
									else
									if((r_sys_run_step==5'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp605[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h9)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==5'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h18)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp374[8:0] );

									end
									else
									if((r_sys_run_step==5'h13)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp470[8:0] );

									end
									else
									if((r_sys_run_step==5'he)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp440[8:0] );

									end
									else
									if((r_sys_run_step==5'h15)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp482[8:0] );

									end
									else
									if((r_sys_run_step==5'h17)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp368[8:0] );

									end
									else
									if((r_sys_run_step==5'h10)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp452[8:0] );

									end
									else
									if((r_sys_run_step==5'h12)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp464[8:0] );

									end
									else
									if((r_sys_run_step==5'h11)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp458[8:0] );

									end
									else
									if((r_sys_run_step==5'h16)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp488[8:0] );

									end
									else
									if((r_sys_run_step==5'h14)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp476[8:0] );

									end
									else
									if((r_sys_run_step==5'hf)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp446[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'he<=r_sys_run_step && r_sys_run_step<=5'h18)) begin
										r_sub00_u_datain <= w_sys_tmp370;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'he<=r_sys_run_step && r_sys_run_step<=5'h18)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp515[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h1: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h2: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								3'h3: begin
									if((r_sys_run_step==5'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((5'h0<=r_sys_run_step && r_sys_run_step<=5'h8)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'ha)) begin
										r_sys_tmp0_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'ha)) begin
										r_sys_tmp0_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h9)) begin
										r_sys_tmp1_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h9)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_tmp2_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h8)) begin
										r_sys_tmp2_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h7)) begin
										r_sys_tmp3_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h7)) begin
										r_sys_tmp3_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_tmp4_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h6)) begin
										r_sys_tmp4_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h5)) begin
										r_sys_tmp5_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h5)) begin
										r_sys_tmp5_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h4)) begin
										r_sys_tmp6_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h4)) begin
										r_sys_tmp6_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3)) begin
										r_sys_tmp7_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h3)) begin
										r_sys_tmp7_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'hb)) begin
										r_sys_tmp8_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								3'h0: begin
									if((r_sys_run_step==5'h2) || (r_sys_run_step==5'hb)) begin
										r_sys_tmp8_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
