/*
TimeStamp:	2016/10/26		15:48
*/


module sub19(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	input  signed  [12:0] i_fld_u_0_addr_0,	
	input          [31:0] i_fld_u_0_datain_0,	
	output         [31:0] o_fld_u_0_dataout_0,	
	input                 i_fld_u_0_r_w_0,	
	input  signed  [12:0] i_fld_result_1_addr_0,	
	input          [31:0] i_fld_result_1_datain_0,	
	output         [31:0] o_fld_result_1_dataout_0,	
	input                 i_fld_result_1_r_w_0	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 1:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 1:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [12:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [12:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [12:0] w_fld_result_1_addr_0;
	wire        [31:0] w_fld_result_1_datain_0;
	wire        [31:0] w_fld_result_1_dataout_0;
	wire               w_fld_result_1_r_w_0;
	wire               w_fld_result_1_ce_0;
	reg  signed [12:0] r_fld_result_1_addr_1;
	reg         [31:0] r_fld_result_1_datain_1;
	wire        [31:0] w_fld_result_1_dataout_1;
	reg                r_fld_result_1_r_w_1;
	wire               w_fld_result_1_ce_1;
	reg  signed [31:0] r_run_k_2;
	reg  signed [31:0] r_run_j_3;
	reg  signed [31:0] r_run_tmpj_4;
	reg         [31:0] r_run_r1_5;
	reg         [31:0] r_run_r2_6;
	reg         [31:0] r_run_dt_7;
	reg         [31:0] r_run_dx_8;
	reg         [31:0] r_run_dy_9;
	reg         [31:0] r_run_q_10;
	reg  signed [31:0] r_run_copy0_j_11;
	reg  signed [31:0] r_run_copy0_j_12;
	reg  signed [31:0] r_run_copy1_j_13;
	reg  signed [31:0] r_run_copy2_j_14;
	reg  signed [31:0] r_run_copy3_j_15;
	reg  signed [31:0] r_run_copy4_j_16;
	reg  signed [31:0] r_run_copy5_j_17;
	reg  signed [31:0] r_run_copy6_j_18;
	reg  signed [31:0] r_run_copy7_j_19;
	reg  signed [31:0] r_run_copy0_j_20;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	wire        [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp4;
	wire signed [31:0] w_sys_tmp6;
	wire               w_sys_tmp7;
	wire               w_sys_tmp8;
	wire signed [31:0] w_sys_tmp9;
	wire signed [31:0] w_sys_tmp12;
	wire signed [31:0] w_sys_tmp13;
	wire        [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire        [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire               w_sys_tmp20;
	wire               w_sys_tmp21;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp26;
	wire signed [31:0] w_sys_tmp27;
	wire        [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp30;
	wire signed [31:0] w_sys_tmp31;
	wire        [31:0] w_sys_tmp34;
	wire signed [31:0] w_sys_tmp35;
	wire signed [31:0] w_sys_tmp36;
	wire signed [31:0] w_sys_tmp102;
	wire               w_sys_tmp103;
	wire               w_sys_tmp104;
	wire signed [31:0] w_sys_tmp105;
	wire signed [31:0] w_sys_tmp106;
	wire signed [31:0] w_sys_tmp107;
	wire               w_sys_tmp108;
	wire               w_sys_tmp109;
	wire signed [31:0] w_sys_tmp110;
	wire signed [31:0] w_sys_tmp113;
	wire signed [31:0] w_sys_tmp114;
	wire signed [31:0] w_sys_tmp115;
	wire        [31:0] w_sys_tmp116;
	wire signed [31:0] w_sys_tmp117;
	wire signed [31:0] w_sys_tmp118;
	wire signed [31:0] w_sys_tmp122;
	wire signed [31:0] w_sys_tmp123;
	wire signed [31:0] w_sys_tmp124;
	wire        [31:0] w_sys_tmp126;
	wire        [31:0] w_sys_tmp127;
	wire        [31:0] w_sys_tmp128;
	wire signed [31:0] w_sys_tmp129;
	wire signed [31:0] w_sys_tmp130;
	wire signed [31:0] w_sys_tmp132;
	wire signed [31:0] w_sys_tmp133;
	wire signed [31:0] w_sys_tmp134;
	wire signed [31:0] w_sys_tmp138;
	wire signed [31:0] w_sys_tmp139;
	wire signed [31:0] w_sys_tmp140;
	wire signed [31:0] w_sys_tmp145;
	wire signed [31:0] w_sys_tmp146;
	wire signed [31:0] w_sys_tmp148;
	wire signed [31:0] w_sys_tmp149;
	wire signed [31:0] w_sys_tmp150;
	wire        [31:0] w_sys_tmp152;
	wire signed [31:0] w_sys_tmp153;
	wire signed [31:0] w_sys_tmp154;
	wire signed [31:0] w_sys_tmp155;
	wire signed [31:0] w_sys_tmp156;
	wire signed [31:0] w_sys_tmp157;
	wire signed [31:0] w_sys_tmp158;
	wire signed [31:0] w_sys_tmp159;
	wire signed [31:0] w_sys_tmp160;
	wire signed [31:0] w_sys_tmp161;
	wire signed [31:0] w_sys_tmp163;
	wire signed [31:0] w_sys_tmp164;
	wire signed [31:0] w_sys_tmp436;
	wire               w_sys_tmp437;
	wire               w_sys_tmp438;
	wire signed [31:0] w_sys_tmp439;
	wire signed [31:0] w_sys_tmp440;
	wire signed [31:0] w_sys_tmp441;
	wire               w_sys_tmp442;
	wire               w_sys_tmp443;
	wire signed [31:0] w_sys_tmp444;
	wire signed [31:0] w_sys_tmp447;
	wire signed [31:0] w_sys_tmp448;
	wire signed [31:0] w_sys_tmp449;
	wire        [31:0] w_sys_tmp450;
	wire signed [31:0] w_sys_tmp451;
	wire signed [31:0] w_sys_tmp452;
	wire signed [31:0] w_sys_tmp454;
	wire signed [31:0] w_sys_tmp455;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 2'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign o_fld_u_0_dataout_0 = w_fld_u_0_dataout_0;
	assign w_fld_u_0_addr_0 = i_fld_u_0_addr_0;
	assign w_fld_u_0_datain_0 = i_fld_u_0_datain_0;
	assign w_fld_u_0_r_w_0 = i_fld_u_0_r_w_0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign o_fld_result_1_dataout_0 = w_fld_result_1_dataout_0;
	assign w_fld_result_1_addr_0 = i_fld_result_1_addr_0;
	assign w_fld_result_1_datain_0 = i_fld_result_1_datain_0;
	assign w_fld_result_1_r_w_0 = i_fld_result_1_r_w_0;
	assign w_fld_result_1_ce_0 = w_sys_ce;
	assign w_fld_result_1_ce_1 = w_sys_ce;
	assign w_sys_tmp1 = 32'h3e4ccccd;
	assign w_sys_tmp3 = 32'h3a03126f;
	assign w_sys_tmp4 = 32'h3d4ccccd;
	assign w_sys_tmp6 = 32'sh00000040;
	assign w_sys_tmp7 = ( !w_sys_tmp8 );
	assign w_sys_tmp8 = (w_sys_tmp9 < r_run_k_2);
	assign w_sys_tmp9 = 32'sh00000061;
	assign w_sys_tmp12 = (w_sys_tmp13 + r_run_k_2);
	assign w_sys_tmp13 = 32'sh00000081;
	assign w_sys_tmp14 = 32'h3f000000;
	assign w_sys_tmp16 = (w_sys_tmp17 + r_run_k_2);
	assign w_sys_tmp17 = 32'sh00004101;
	assign w_sys_tmp18 = 32'h0;
	assign w_sys_tmp19 = (r_run_k_2 + w_sys_intOne);
	assign w_sys_tmp20 = ( !w_sys_tmp21 );
	assign w_sys_tmp21 = (w_sys_tmp22 < r_run_j_3);
	assign w_sys_tmp22 = 32'sh00000012;
	assign w_sys_tmp25 = (w_sys_tmp26 + w_sys_intOne);
	assign w_sys_tmp26 = (r_run_j_3 * w_sys_tmp27);
	assign w_sys_tmp27 = 32'sh00000081;
	assign w_sys_tmp28 = 32'h3f800000;
	assign w_sys_tmp30 = (w_sys_tmp31 + w_sys_tmp27);
	assign w_sys_tmp31 = (r_run_copy0_j_11 * w_sys_tmp27);
	assign w_sys_tmp34 = 32'h0;
	assign w_sys_tmp35 = (r_run_copy0_j_11 + w_sys_intOne);
	assign w_sys_tmp36 = (r_run_j_3 + w_sys_intOne);
	assign w_sys_tmp102 = 32'sh00000041;
	assign w_sys_tmp103 = ( !w_sys_tmp104 );
	assign w_sys_tmp104 = (w_sys_tmp105 < r_run_k_2);
	assign w_sys_tmp105 = 32'sh00000060;
	assign w_sys_tmp106 = (r_run_k_2 + w_sys_intOne);
	assign w_sys_tmp107 = 32'sh00000002;
	assign w_sys_tmp108 = ( !w_sys_tmp109 );
	assign w_sys_tmp109 = (w_sys_tmp110 < r_run_j_3);
	assign w_sys_tmp110 = 32'sh00000011;
	assign w_sys_tmp113 = (w_sys_tmp114 + r_run_k_2);
	assign w_sys_tmp114 = (r_run_j_3 * w_sys_tmp115);
	assign w_sys_tmp115 = 32'sh00000081;
	assign w_sys_tmp116 = w_ip_AddFloat_result_0;
	assign w_sys_tmp117 = (w_sys_tmp118 + r_run_k_2);
	assign w_sys_tmp118 = (r_run_copy7_j_19 * w_sys_tmp115);
	assign w_sys_tmp122 = (w_sys_tmp123 + r_run_k_2);
	assign w_sys_tmp123 = (w_sys_tmp124 * w_sys_tmp115);
	assign w_sys_tmp124 = (r_run_copy6_j_18 + w_sys_intOne);
	assign w_sys_tmp126 = w_ip_MultFloat_product_0;
	assign w_sys_tmp127 = 32'h40000000;
	assign w_sys_tmp128 = w_fld_u_0_dataout_1;
	assign w_sys_tmp129 = (w_sys_tmp130 + r_run_k_2);
	assign w_sys_tmp130 = (r_run_copy5_j_17 * w_sys_tmp115);
	assign w_sys_tmp132 = (w_sys_tmp133 + r_run_k_2);
	assign w_sys_tmp133 = (w_sys_tmp134 * w_sys_tmp115);
	assign w_sys_tmp134 = (r_run_copy4_j_16 - w_sys_intOne);
	assign w_sys_tmp138 = (w_sys_tmp139 + w_sys_intOne);
	assign w_sys_tmp139 = (w_sys_tmp140 + r_run_k_2);
	assign w_sys_tmp140 = (r_run_copy3_j_15 * w_sys_tmp115);
	assign w_sys_tmp145 = (w_sys_tmp146 + r_run_k_2);
	assign w_sys_tmp146 = (r_run_copy2_j_14 * w_sys_tmp115);
	assign w_sys_tmp148 = (w_sys_tmp149 - w_sys_intOne);
	assign w_sys_tmp149 = (w_sys_tmp150 + r_run_k_2);
	assign w_sys_tmp150 = (r_run_copy1_j_13 * w_sys_tmp115);
	assign w_sys_tmp152 = 32'h42c80000;
	assign w_sys_tmp153 = (r_run_copy0_j_12 + w_sys_tmp154);
	assign w_sys_tmp154 = 32'sh0000006e;
	assign w_sys_tmp155 = (r_run_k_2 - w_sys_intOne);
	assign w_sys_tmp156 = (r_run_copy0_j_12 + w_sys_intOne);
	assign w_sys_tmp157 = (r_run_copy1_j_13 + w_sys_intOne);
	assign w_sys_tmp158 = (r_run_copy2_j_14 + w_sys_intOne);
	assign w_sys_tmp159 = (r_run_copy3_j_15 + w_sys_intOne);
	assign w_sys_tmp160 = (r_run_copy4_j_16 + w_sys_intOne);
	assign w_sys_tmp161 = (r_run_copy5_j_17 + w_sys_intOne);
	assign w_sys_tmp163 = (r_run_copy7_j_19 + w_sys_intOne);
	assign w_sys_tmp164 = (r_run_j_3 + w_sys_intOne);
	assign w_sys_tmp436 = 32'sh00000041;
	assign w_sys_tmp437 = ( !w_sys_tmp438 );
	assign w_sys_tmp438 = (w_sys_tmp439 < r_run_k_2);
	assign w_sys_tmp439 = 32'sh00000060;
	assign w_sys_tmp440 = (r_run_k_2 + w_sys_intOne);
	assign w_sys_tmp441 = 32'sh00000002;
	assign w_sys_tmp442 = ( !w_sys_tmp443 );
	assign w_sys_tmp443 = (w_sys_tmp444 < r_run_j_3);
	assign w_sys_tmp444 = 32'sh00000011;
	assign w_sys_tmp447 = (w_sys_tmp448 + r_run_k_2);
	assign w_sys_tmp448 = (r_run_j_3 * w_sys_tmp449);
	assign w_sys_tmp449 = 32'sh00000081;
	assign w_sys_tmp450 = w_fld_result_1_dataout_1;
	assign w_sys_tmp451 = (w_sys_tmp452 + r_run_k_2);
	assign w_sys_tmp452 = (r_run_copy0_j_20 * w_sys_tmp449);
	assign w_sys_tmp454 = (r_run_copy0_j_20 + w_sys_intOne);
	assign w_sys_tmp455 = (r_run_j_3 + w_sys_intOne);


	DualPortRAM #(.DWIDTH(32), .AWIDTH(13), .WORDS(4515) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(13), .WORDS(4515) )
		dpram_result_1(
			.clk (clock),
			.ce_0 (w_fld_result_1_ce_0),
			.addr_0 (w_fld_result_1_addr_0),
			.datain_0 (w_fld_result_1_datain_0),
			.dataout_0 (w_fld_result_1_dataout_0),
			.r_w_0 (w_fld_result_1_r_w_0),
			.ce_1 (w_fld_result_1_ce_1),
			.addr_1 (r_fld_result_1_addr_1),
			.datain_1 (r_fld_result_1_datain_1),
			.dataout_1 (w_fld_result_1_dataout_1),
			.r_w_1 (r_fld_result_1_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1e) || (r_sys_run_step==7'h35)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h13) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h36)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2f)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h45)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp116;

									end
									else
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h3b)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h29) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h37)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h27)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h17) || (r_sys_run_step==7'h2e)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h22) || (r_sys_run_step==7'h32)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h20)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp14_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h18)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h1c) || (r_sys_run_step==7'h26)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'h15) || (r_sys_run_step==7'h1f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h27) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'h22) || (r_sys_run_step==7'h3b)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp126;

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'h20) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h40)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==7'h19) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h45)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'h23) || (r_sys_run_step==7'h2d)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
									else
									if((r_sys_run_step==7'h2a) || (r_sys_run_step==7'h34)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp126[31], w_sys_tmp126[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h6)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dt_7;

									end
									else
									if((r_sys_run_step==7'h1b) || (r_sys_run_step==7'h26)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h1d) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h39)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r2_6;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2d)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==7'h8) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h33)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2e)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'h13) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h36)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r1_5;

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2a)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp127;

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h29) || (r_sys_run_step==7'h30)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp152;

									end
									else
									if((r_sys_run_step==7'h8) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_dx_8;

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h30)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h29)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_dy_9;

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2a)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp128;

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'h11) || (r_sys_run_step==7'h31)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'h13) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h39)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp116;

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h1f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp153;

									end
									else
									if((7'h6<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp155;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h26: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7) ? 6'h8 : 6'ha);

									end
								end

							endcase
						end

						6'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'hb;

									end
								end

							endcase
						end

						6'hb: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp20) ? 6'he : 6'h10);

									end
								end

							endcase
						end

						6'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_run_phase <= 6'hb;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h11;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp103) ? 6'h15 : 6'h1b);

									end
								end

							endcase
						end

						6'h12: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h11;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h16;

									end
								end

							endcase
						end

						6'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp108) ? 6'h19 : 6'h12);

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h4a)) begin
										r_sys_run_phase <= 6'h16;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h1c;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp437) ? 6'h20 : 6'h26);

									end
								end

							endcase
						end

						6'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h1c;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp442) ? 6'h24 : 6'h1d);

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h26: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'hb: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h12: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h4a)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'hb: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'ha)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h12: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h4a)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h49)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h26: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp16[12:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp12[12:0] );

									end
								end

							endcase
						end

						6'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h2) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp25[12:0] );

									end
									else
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp30[12:0] );

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp148[12:0] );

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp138[12:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp132[12:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp145[12:0] );

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp129[12:0] );

									end
									else
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp122[12:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp117[12:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp447[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp18;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp14;

									end
								end

							endcase
						end

						6'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h2) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'ha)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp28;

									end
									else
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp34;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp450;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h29)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h26: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_result_1_addr_1 <= 13'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h4a)) begin
										r_fld_result_1_addr_1 <= $signed( w_sys_tmp113[12:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_fld_result_1_addr_1 <= $signed( w_sys_tmp451[12:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h4a)) begin
										r_fld_result_1_datain_1 <= w_sys_tmp116;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_result_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h4a)) begin
										r_fld_result_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_fld_result_1_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h26: begin
							r_fld_result_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_2 <= w_sys_tmp6;

									end
								end

							endcase
						end

						6'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_run_k_2 <= w_sys_tmp19;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_2 <= w_sys_tmp102;

									end
								end

							endcase
						end

						6'h12: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_2 <= w_sys_tmp106;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_2 <= w_sys_tmp436;

									end
								end

							endcase
						end

						6'h1d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_2 <= w_sys_tmp440;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_3 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h2) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'ha)) begin
										r_run_j_3 <= w_sys_tmp36;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_3 <= w_sys_tmp107;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h4a)) begin
										r_run_j_3 <= w_sys_tmp164;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_3 <= w_sys_tmp441;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_run_j_3 <= w_sys_tmp455;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r1_5 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r2_6 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dt_7 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dx_8 <= w_sys_tmp4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dy_9 <= w_sys_tmp4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'ha: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_11 <= r_run_j_3;

									end
								end

							endcase
						end

						6'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb)) begin
										r_run_copy0_j_11 <= w_sys_tmp35;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_12 <= r_run_j_3;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_run_copy0_j_12 <= w_sys_tmp156;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_13 <= r_run_j_3;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h29)) begin
										r_run_copy1_j_13 <= w_sys_tmp157;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_14 <= r_run_j_3;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h28)) begin
										r_run_copy2_j_14 <= w_sys_tmp158;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_15 <= r_run_j_3;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h27)) begin
										r_run_copy3_j_15 <= w_sys_tmp159;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_16 <= r_run_j_3;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h26)) begin
										r_run_copy4_j_16 <= w_sys_tmp160;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy5_j_17 <= r_run_j_3;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h25)) begin
										r_run_copy5_j_17 <= w_sys_tmp161;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy6_j_18 <= r_run_j_3;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h24)) begin
										r_run_copy6_j_18 <= w_sys_tmp124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy7_j_19 <= r_run_j_3;

									end
								end

							endcase
						end

						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h23)) begin
										r_run_copy7_j_19 <= w_sys_tmp163;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h20: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_20 <= r_run_j_3;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_run_copy0_j_20 <= w_sys_tmp454;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h12)) begin
										r_sys_tmp0_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hf)) begin
										r_sys_tmp1_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'he)) begin
										r_sys_tmp2_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_tmp3_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h8) || (r_sys_run_step==7'h11)) begin
										r_sys_tmp5_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'h10)) begin
										r_sys_tmp6_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h15) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29)) begin
										r_sys_tmp7_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h28)) begin
										r_sys_tmp8_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h8) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h17)) begin
										r_sys_tmp9_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h24)) begin
										r_sys_tmp10_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h24) || (r_sys_run_step==7'h2b)) begin
										r_sys_tmp11_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sys_tmp11_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1e) || (r_sys_run_step==7'h27)) begin
										r_sys_tmp12_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp12_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1e)) begin
										r_sys_tmp13_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h2b)) begin
										r_sys_tmp14_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h25)) begin
										r_sys_tmp15_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp16_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==7'h14) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h29)) begin
										r_sys_tmp16_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h2e)) begin
										r_sys_tmp17_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h26)) begin
										r_sys_tmp17_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h35)) begin
										r_sys_tmp18_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp18_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h36)) begin
										r_sys_tmp19_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h38)) begin
										r_sys_tmp20_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h3e)) begin
										r_sys_tmp21_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
