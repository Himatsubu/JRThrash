/*
TimeStamp:	2016/5/18		3:32
*/


module P3_2dim(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg  signed [31:0] r_ip_DivInt_dividend_0;
	reg  signed [31:0] r_ip_DivInt_divisor_0;
	wire signed [31:0] w_ip_DivInt_quotient_0;
	wire signed [31:0] w_ip_DivInt_fractional_0;
	reg  signed [31:0] r_ip_DivInt_dividend_1;
	reg  signed [31:0] r_ip_DivInt_divisor_1;
	wire signed [31:0] w_ip_DivInt_quotient_1;
	wire signed [31:0] w_ip_DivInt_fractional_1;
	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 7:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 7:0] w_sys_run_step_p1;
	wire signed [ 9:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [ 9:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [ 9:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [ 9:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [ 9:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [ 9:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [ 9:0] w_fld_V_3_addr_0;
	wire        [31:0] w_fld_V_3_datain_0;
	wire        [31:0] w_fld_V_3_dataout_0;
	wire               w_fld_V_3_r_w_0;
	wire               w_fld_V_3_ce_0;
	reg  signed [ 9:0] r_fld_V_3_addr_1;
	reg         [31:0] r_fld_V_3_datain_1;
	wire        [31:0] w_fld_V_3_dataout_1;
	reg                r_fld_V_3_r_w_1;
	wire               w_fld_V_3_ce_1;
	reg  signed [31:0] r_run_k_29;
	reg  signed [31:0] r_run_j_30;
	reg  signed [31:0] r_run_n_31;
	reg  signed [31:0] r_run_mx_32;
	reg  signed [31:0] r_run_my_33;
	reg         [31:0] r_run_dt_34;
	reg         [31:0] r_run_dx_35;
	reg         [31:0] r_run_dy_36;
	reg         [31:0] r_run_r1_37;
	reg         [31:0] r_run_r2_38;
	reg         [31:0] r_run_r3_39;
	reg         [31:0] r_run_r4_40;
	reg         [31:0] r_run_YY_41;
	reg  signed [31:0] r_run_kx_42;
	reg  signed [31:0] r_run_ky_43;
	reg  signed [31:0] r_run_nlast_44;
	reg  signed [31:0] r_run_copy0_j_45;
	reg  signed [31:0] r_run_copy1_j_46;
	reg  signed [31:0] r_run_copy2_j_47;
	reg  signed [31:0] r_run_copy0_j_48;
	reg                r_sub19_run_req;
	wire               w_sub19_run_busy;
	wire signed [ 9:0] w_sub19_T_addr;
	reg  signed [ 9:0] r_sub19_T_addr;
	wire        [31:0] w_sub19_T_datain;
	reg         [31:0] r_sub19_T_datain;
	wire        [31:0] w_sub19_T_dataout;
	wire               w_sub19_T_r_w;
	reg                r_sub19_T_r_w;
	wire signed [ 9:0] w_sub19_V_addr;
	reg  signed [ 9:0] r_sub19_V_addr;
	wire        [31:0] w_sub19_V_datain;
	reg         [31:0] r_sub19_V_datain;
	wire        [31:0] w_sub19_V_dataout;
	wire               w_sub19_V_r_w;
	reg                r_sub19_V_r_w;
	wire signed [ 9:0] w_sub19_U_addr;
	reg  signed [ 9:0] r_sub19_U_addr;
	wire        [31:0] w_sub19_U_datain;
	reg         [31:0] r_sub19_U_datain;
	wire        [31:0] w_sub19_U_dataout;
	wire               w_sub19_U_r_w;
	reg                r_sub19_U_r_w;
	wire signed [ 9:0] w_sub19_result_addr;
	reg  signed [ 9:0] r_sub19_result_addr;
	wire        [31:0] w_sub19_result_datain;
	reg         [31:0] r_sub19_result_datain;
	wire        [31:0] w_sub19_result_dataout;
	wire               w_sub19_result_r_w;
	reg                r_sub19_result_r_w;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [ 9:0] w_sub09_T_addr;
	reg  signed [ 9:0] r_sub09_T_addr;
	wire        [31:0] w_sub09_T_datain;
	reg         [31:0] r_sub09_T_datain;
	wire        [31:0] w_sub09_T_dataout;
	wire               w_sub09_T_r_w;
	reg                r_sub09_T_r_w;
	wire signed [ 9:0] w_sub09_V_addr;
	reg  signed [ 9:0] r_sub09_V_addr;
	wire        [31:0] w_sub09_V_datain;
	reg         [31:0] r_sub09_V_datain;
	wire        [31:0] w_sub09_V_dataout;
	wire               w_sub09_V_r_w;
	reg                r_sub09_V_r_w;
	wire signed [ 9:0] w_sub09_U_addr;
	reg  signed [ 9:0] r_sub09_U_addr;
	wire        [31:0] w_sub09_U_datain;
	reg         [31:0] r_sub09_U_datain;
	wire        [31:0] w_sub09_U_dataout;
	wire               w_sub09_U_r_w;
	reg                r_sub09_U_r_w;
	wire signed [ 9:0] w_sub09_result_addr;
	reg  signed [ 9:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [ 9:0] w_sub08_T_addr;
	reg  signed [ 9:0] r_sub08_T_addr;
	wire        [31:0] w_sub08_T_datain;
	reg         [31:0] r_sub08_T_datain;
	wire        [31:0] w_sub08_T_dataout;
	wire               w_sub08_T_r_w;
	reg                r_sub08_T_r_w;
	wire signed [ 9:0] w_sub08_V_addr;
	reg  signed [ 9:0] r_sub08_V_addr;
	wire        [31:0] w_sub08_V_datain;
	reg         [31:0] r_sub08_V_datain;
	wire        [31:0] w_sub08_V_dataout;
	wire               w_sub08_V_r_w;
	reg                r_sub08_V_r_w;
	wire signed [ 9:0] w_sub08_U_addr;
	reg  signed [ 9:0] r_sub08_U_addr;
	wire        [31:0] w_sub08_U_datain;
	reg         [31:0] r_sub08_U_datain;
	wire        [31:0] w_sub08_U_dataout;
	wire               w_sub08_U_r_w;
	reg                r_sub08_U_r_w;
	wire signed [ 9:0] w_sub08_result_addr;
	reg  signed [ 9:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub24_run_req;
	wire               w_sub24_run_busy;
	wire signed [ 9:0] w_sub24_T_addr;
	reg  signed [ 9:0] r_sub24_T_addr;
	wire        [31:0] w_sub24_T_datain;
	reg         [31:0] r_sub24_T_datain;
	wire        [31:0] w_sub24_T_dataout;
	wire               w_sub24_T_r_w;
	reg                r_sub24_T_r_w;
	wire signed [ 9:0] w_sub24_V_addr;
	reg  signed [ 9:0] r_sub24_V_addr;
	wire        [31:0] w_sub24_V_datain;
	reg         [31:0] r_sub24_V_datain;
	wire        [31:0] w_sub24_V_dataout;
	wire               w_sub24_V_r_w;
	reg                r_sub24_V_r_w;
	wire signed [ 9:0] w_sub24_U_addr;
	reg  signed [ 9:0] r_sub24_U_addr;
	wire        [31:0] w_sub24_U_datain;
	reg         [31:0] r_sub24_U_datain;
	wire        [31:0] w_sub24_U_dataout;
	wire               w_sub24_U_r_w;
	reg                r_sub24_U_r_w;
	wire signed [ 9:0] w_sub24_result_addr;
	reg  signed [ 9:0] r_sub24_result_addr;
	wire        [31:0] w_sub24_result_datain;
	reg         [31:0] r_sub24_result_datain;
	wire        [31:0] w_sub24_result_dataout;
	wire               w_sub24_result_r_w;
	reg                r_sub24_result_r_w;
	reg                r_sub22_run_req;
	wire               w_sub22_run_busy;
	wire signed [ 9:0] w_sub22_T_addr;
	reg  signed [ 9:0] r_sub22_T_addr;
	wire        [31:0] w_sub22_T_datain;
	reg         [31:0] r_sub22_T_datain;
	wire        [31:0] w_sub22_T_dataout;
	wire               w_sub22_T_r_w;
	reg                r_sub22_T_r_w;
	wire signed [ 9:0] w_sub22_V_addr;
	reg  signed [ 9:0] r_sub22_V_addr;
	wire        [31:0] w_sub22_V_datain;
	reg         [31:0] r_sub22_V_datain;
	wire        [31:0] w_sub22_V_dataout;
	wire               w_sub22_V_r_w;
	reg                r_sub22_V_r_w;
	wire signed [ 9:0] w_sub22_U_addr;
	reg  signed [ 9:0] r_sub22_U_addr;
	wire        [31:0] w_sub22_U_datain;
	reg         [31:0] r_sub22_U_datain;
	wire        [31:0] w_sub22_U_dataout;
	wire               w_sub22_U_r_w;
	reg                r_sub22_U_r_w;
	wire signed [ 9:0] w_sub22_result_addr;
	reg  signed [ 9:0] r_sub22_result_addr;
	wire        [31:0] w_sub22_result_datain;
	reg         [31:0] r_sub22_result_datain;
	wire        [31:0] w_sub22_result_dataout;
	wire               w_sub22_result_r_w;
	reg                r_sub22_result_r_w;
	reg                r_sub23_run_req;
	wire               w_sub23_run_busy;
	wire signed [ 9:0] w_sub23_T_addr;
	reg  signed [ 9:0] r_sub23_T_addr;
	wire        [31:0] w_sub23_T_datain;
	reg         [31:0] r_sub23_T_datain;
	wire        [31:0] w_sub23_T_dataout;
	wire               w_sub23_T_r_w;
	reg                r_sub23_T_r_w;
	wire signed [ 9:0] w_sub23_V_addr;
	reg  signed [ 9:0] r_sub23_V_addr;
	wire        [31:0] w_sub23_V_datain;
	reg         [31:0] r_sub23_V_datain;
	wire        [31:0] w_sub23_V_dataout;
	wire               w_sub23_V_r_w;
	reg                r_sub23_V_r_w;
	wire signed [ 9:0] w_sub23_U_addr;
	reg  signed [ 9:0] r_sub23_U_addr;
	wire        [31:0] w_sub23_U_datain;
	reg         [31:0] r_sub23_U_datain;
	wire        [31:0] w_sub23_U_dataout;
	wire               w_sub23_U_r_w;
	reg                r_sub23_U_r_w;
	wire signed [ 9:0] w_sub23_result_addr;
	reg  signed [ 9:0] r_sub23_result_addr;
	wire        [31:0] w_sub23_result_datain;
	reg         [31:0] r_sub23_result_datain;
	wire        [31:0] w_sub23_result_dataout;
	wire               w_sub23_result_r_w;
	reg                r_sub23_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [ 9:0] w_sub12_T_addr;
	reg  signed [ 9:0] r_sub12_T_addr;
	wire        [31:0] w_sub12_T_datain;
	reg         [31:0] r_sub12_T_datain;
	wire        [31:0] w_sub12_T_dataout;
	wire               w_sub12_T_r_w;
	reg                r_sub12_T_r_w;
	wire signed [ 9:0] w_sub12_V_addr;
	reg  signed [ 9:0] r_sub12_V_addr;
	wire        [31:0] w_sub12_V_datain;
	reg         [31:0] r_sub12_V_datain;
	wire        [31:0] w_sub12_V_dataout;
	wire               w_sub12_V_r_w;
	reg                r_sub12_V_r_w;
	wire signed [ 9:0] w_sub12_U_addr;
	reg  signed [ 9:0] r_sub12_U_addr;
	wire        [31:0] w_sub12_U_datain;
	reg         [31:0] r_sub12_U_datain;
	wire        [31:0] w_sub12_U_dataout;
	wire               w_sub12_U_r_w;
	reg                r_sub12_U_r_w;
	wire signed [ 9:0] w_sub12_result_addr;
	reg  signed [ 9:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 9:0] w_sub03_T_addr;
	reg  signed [ 9:0] r_sub03_T_addr;
	wire        [31:0] w_sub03_T_datain;
	reg         [31:0] r_sub03_T_datain;
	wire        [31:0] w_sub03_T_dataout;
	wire               w_sub03_T_r_w;
	reg                r_sub03_T_r_w;
	wire signed [ 9:0] w_sub03_V_addr;
	reg  signed [ 9:0] r_sub03_V_addr;
	wire        [31:0] w_sub03_V_datain;
	reg         [31:0] r_sub03_V_datain;
	wire        [31:0] w_sub03_V_dataout;
	wire               w_sub03_V_r_w;
	reg                r_sub03_V_r_w;
	wire signed [ 9:0] w_sub03_U_addr;
	reg  signed [ 9:0] r_sub03_U_addr;
	wire        [31:0] w_sub03_U_datain;
	reg         [31:0] r_sub03_U_datain;
	wire        [31:0] w_sub03_U_dataout;
	wire               w_sub03_U_r_w;
	reg                r_sub03_U_r_w;
	wire signed [ 9:0] w_sub03_result_addr;
	reg  signed [ 9:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 9:0] w_sub02_T_addr;
	reg  signed [ 9:0] r_sub02_T_addr;
	wire        [31:0] w_sub02_T_datain;
	reg         [31:0] r_sub02_T_datain;
	wire        [31:0] w_sub02_T_dataout;
	wire               w_sub02_T_r_w;
	reg                r_sub02_T_r_w;
	wire signed [ 9:0] w_sub02_V_addr;
	reg  signed [ 9:0] r_sub02_V_addr;
	wire        [31:0] w_sub02_V_datain;
	reg         [31:0] r_sub02_V_datain;
	wire        [31:0] w_sub02_V_dataout;
	wire               w_sub02_V_r_w;
	reg                r_sub02_V_r_w;
	wire signed [ 9:0] w_sub02_U_addr;
	reg  signed [ 9:0] r_sub02_U_addr;
	wire        [31:0] w_sub02_U_datain;
	reg         [31:0] r_sub02_U_datain;
	wire        [31:0] w_sub02_U_dataout;
	wire               w_sub02_U_r_w;
	reg                r_sub02_U_r_w;
	wire signed [ 9:0] w_sub02_result_addr;
	reg  signed [ 9:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [ 9:0] w_sub11_T_addr;
	reg  signed [ 9:0] r_sub11_T_addr;
	wire        [31:0] w_sub11_T_datain;
	reg         [31:0] r_sub11_T_datain;
	wire        [31:0] w_sub11_T_dataout;
	wire               w_sub11_T_r_w;
	reg                r_sub11_T_r_w;
	wire signed [ 9:0] w_sub11_V_addr;
	reg  signed [ 9:0] r_sub11_V_addr;
	wire        [31:0] w_sub11_V_datain;
	reg         [31:0] r_sub11_V_datain;
	wire        [31:0] w_sub11_V_dataout;
	wire               w_sub11_V_r_w;
	reg                r_sub11_V_r_w;
	wire signed [ 9:0] w_sub11_U_addr;
	reg  signed [ 9:0] r_sub11_U_addr;
	wire        [31:0] w_sub11_U_datain;
	reg         [31:0] r_sub11_U_datain;
	wire        [31:0] w_sub11_U_dataout;
	wire               w_sub11_U_r_w;
	reg                r_sub11_U_r_w;
	wire signed [ 9:0] w_sub11_result_addr;
	reg  signed [ 9:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [ 9:0] w_sub14_T_addr;
	reg  signed [ 9:0] r_sub14_T_addr;
	wire        [31:0] w_sub14_T_datain;
	reg         [31:0] r_sub14_T_datain;
	wire        [31:0] w_sub14_T_dataout;
	wire               w_sub14_T_r_w;
	reg                r_sub14_T_r_w;
	wire signed [ 9:0] w_sub14_V_addr;
	reg  signed [ 9:0] r_sub14_V_addr;
	wire        [31:0] w_sub14_V_datain;
	reg         [31:0] r_sub14_V_datain;
	wire        [31:0] w_sub14_V_dataout;
	wire               w_sub14_V_r_w;
	reg                r_sub14_V_r_w;
	wire signed [ 9:0] w_sub14_U_addr;
	reg  signed [ 9:0] r_sub14_U_addr;
	wire        [31:0] w_sub14_U_datain;
	reg         [31:0] r_sub14_U_datain;
	wire        [31:0] w_sub14_U_dataout;
	wire               w_sub14_U_r_w;
	reg                r_sub14_U_r_w;
	wire signed [ 9:0] w_sub14_result_addr;
	reg  signed [ 9:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 9:0] w_sub01_T_addr;
	reg  signed [ 9:0] r_sub01_T_addr;
	wire        [31:0] w_sub01_T_datain;
	reg         [31:0] r_sub01_T_datain;
	wire        [31:0] w_sub01_T_dataout;
	wire               w_sub01_T_r_w;
	reg                r_sub01_T_r_w;
	wire signed [ 9:0] w_sub01_V_addr;
	reg  signed [ 9:0] r_sub01_V_addr;
	wire        [31:0] w_sub01_V_datain;
	reg         [31:0] r_sub01_V_datain;
	wire        [31:0] w_sub01_V_dataout;
	wire               w_sub01_V_r_w;
	reg                r_sub01_V_r_w;
	wire signed [ 9:0] w_sub01_U_addr;
	reg  signed [ 9:0] r_sub01_U_addr;
	wire        [31:0] w_sub01_U_datain;
	reg         [31:0] r_sub01_U_datain;
	wire        [31:0] w_sub01_U_dataout;
	wire               w_sub01_U_r_w;
	reg                r_sub01_U_r_w;
	wire signed [ 9:0] w_sub01_result_addr;
	reg  signed [ 9:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 9:0] w_sub00_T_addr;
	reg  signed [ 9:0] r_sub00_T_addr;
	wire        [31:0] w_sub00_T_datain;
	reg         [31:0] r_sub00_T_datain;
	wire        [31:0] w_sub00_T_dataout;
	wire               w_sub00_T_r_w;
	reg                r_sub00_T_r_w;
	wire signed [ 9:0] w_sub00_V_addr;
	reg  signed [ 9:0] r_sub00_V_addr;
	wire        [31:0] w_sub00_V_datain;
	reg         [31:0] r_sub00_V_datain;
	wire        [31:0] w_sub00_V_dataout;
	wire               w_sub00_V_r_w;
	reg                r_sub00_V_r_w;
	wire signed [ 9:0] w_sub00_U_addr;
	reg  signed [ 9:0] r_sub00_U_addr;
	wire        [31:0] w_sub00_U_datain;
	reg         [31:0] r_sub00_U_datain;
	wire        [31:0] w_sub00_U_dataout;
	wire               w_sub00_U_r_w;
	reg                r_sub00_U_r_w;
	wire signed [ 9:0] w_sub00_result_addr;
	reg  signed [ 9:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [ 9:0] w_sub13_T_addr;
	reg  signed [ 9:0] r_sub13_T_addr;
	wire        [31:0] w_sub13_T_datain;
	reg         [31:0] r_sub13_T_datain;
	wire        [31:0] w_sub13_T_dataout;
	wire               w_sub13_T_r_w;
	reg                r_sub13_T_r_w;
	wire signed [ 9:0] w_sub13_V_addr;
	reg  signed [ 9:0] r_sub13_V_addr;
	wire        [31:0] w_sub13_V_datain;
	reg         [31:0] r_sub13_V_datain;
	wire        [31:0] w_sub13_V_dataout;
	wire               w_sub13_V_r_w;
	reg                r_sub13_V_r_w;
	wire signed [ 9:0] w_sub13_U_addr;
	reg  signed [ 9:0] r_sub13_U_addr;
	wire        [31:0] w_sub13_U_datain;
	reg         [31:0] r_sub13_U_datain;
	wire        [31:0] w_sub13_U_dataout;
	wire               w_sub13_U_r_w;
	reg                r_sub13_U_r_w;
	wire signed [ 9:0] w_sub13_result_addr;
	reg  signed [ 9:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [ 9:0] w_sub07_T_addr;
	reg  signed [ 9:0] r_sub07_T_addr;
	wire        [31:0] w_sub07_T_datain;
	reg         [31:0] r_sub07_T_datain;
	wire        [31:0] w_sub07_T_dataout;
	wire               w_sub07_T_r_w;
	reg                r_sub07_T_r_w;
	wire signed [ 9:0] w_sub07_V_addr;
	reg  signed [ 9:0] r_sub07_V_addr;
	wire        [31:0] w_sub07_V_datain;
	reg         [31:0] r_sub07_V_datain;
	wire        [31:0] w_sub07_V_dataout;
	wire               w_sub07_V_r_w;
	reg                r_sub07_V_r_w;
	wire signed [ 9:0] w_sub07_U_addr;
	reg  signed [ 9:0] r_sub07_U_addr;
	wire        [31:0] w_sub07_U_datain;
	reg         [31:0] r_sub07_U_datain;
	wire        [31:0] w_sub07_U_dataout;
	wire               w_sub07_U_r_w;
	reg                r_sub07_U_r_w;
	wire signed [ 9:0] w_sub07_result_addr;
	reg  signed [ 9:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub16_run_req;
	wire               w_sub16_run_busy;
	wire signed [ 9:0] w_sub16_T_addr;
	reg  signed [ 9:0] r_sub16_T_addr;
	wire        [31:0] w_sub16_T_datain;
	reg         [31:0] r_sub16_T_datain;
	wire        [31:0] w_sub16_T_dataout;
	wire               w_sub16_T_r_w;
	reg                r_sub16_T_r_w;
	wire signed [ 9:0] w_sub16_V_addr;
	reg  signed [ 9:0] r_sub16_V_addr;
	wire        [31:0] w_sub16_V_datain;
	reg         [31:0] r_sub16_V_datain;
	wire        [31:0] w_sub16_V_dataout;
	wire               w_sub16_V_r_w;
	reg                r_sub16_V_r_w;
	wire signed [ 9:0] w_sub16_U_addr;
	reg  signed [ 9:0] r_sub16_U_addr;
	wire        [31:0] w_sub16_U_datain;
	reg         [31:0] r_sub16_U_datain;
	wire        [31:0] w_sub16_U_dataout;
	wire               w_sub16_U_r_w;
	reg                r_sub16_U_r_w;
	wire signed [ 9:0] w_sub16_result_addr;
	reg  signed [ 9:0] r_sub16_result_addr;
	wire        [31:0] w_sub16_result_datain;
	reg         [31:0] r_sub16_result_datain;
	wire        [31:0] w_sub16_result_dataout;
	wire               w_sub16_result_r_w;
	reg                r_sub16_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [ 9:0] w_sub06_T_addr;
	reg  signed [ 9:0] r_sub06_T_addr;
	wire        [31:0] w_sub06_T_datain;
	reg         [31:0] r_sub06_T_datain;
	wire        [31:0] w_sub06_T_dataout;
	wire               w_sub06_T_r_w;
	reg                r_sub06_T_r_w;
	wire signed [ 9:0] w_sub06_V_addr;
	reg  signed [ 9:0] r_sub06_V_addr;
	wire        [31:0] w_sub06_V_datain;
	reg         [31:0] r_sub06_V_datain;
	wire        [31:0] w_sub06_V_dataout;
	wire               w_sub06_V_r_w;
	reg                r_sub06_V_r_w;
	wire signed [ 9:0] w_sub06_U_addr;
	reg  signed [ 9:0] r_sub06_U_addr;
	wire        [31:0] w_sub06_U_datain;
	reg         [31:0] r_sub06_U_datain;
	wire        [31:0] w_sub06_U_dataout;
	wire               w_sub06_U_r_w;
	reg                r_sub06_U_r_w;
	wire signed [ 9:0] w_sub06_result_addr;
	reg  signed [ 9:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [ 9:0] w_sub15_T_addr;
	reg  signed [ 9:0] r_sub15_T_addr;
	wire        [31:0] w_sub15_T_datain;
	reg         [31:0] r_sub15_T_datain;
	wire        [31:0] w_sub15_T_dataout;
	wire               w_sub15_T_r_w;
	reg                r_sub15_T_r_w;
	wire signed [ 9:0] w_sub15_V_addr;
	reg  signed [ 9:0] r_sub15_V_addr;
	wire        [31:0] w_sub15_V_datain;
	reg         [31:0] r_sub15_V_datain;
	wire        [31:0] w_sub15_V_dataout;
	wire               w_sub15_V_r_w;
	reg                r_sub15_V_r_w;
	wire signed [ 9:0] w_sub15_U_addr;
	reg  signed [ 9:0] r_sub15_U_addr;
	wire        [31:0] w_sub15_U_datain;
	reg         [31:0] r_sub15_U_datain;
	wire        [31:0] w_sub15_U_dataout;
	wire               w_sub15_U_r_w;
	reg                r_sub15_U_r_w;
	wire signed [ 9:0] w_sub15_result_addr;
	reg  signed [ 9:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [ 9:0] w_sub05_T_addr;
	reg  signed [ 9:0] r_sub05_T_addr;
	wire        [31:0] w_sub05_T_datain;
	reg         [31:0] r_sub05_T_datain;
	wire        [31:0] w_sub05_T_dataout;
	wire               w_sub05_T_r_w;
	reg                r_sub05_T_r_w;
	wire signed [ 9:0] w_sub05_V_addr;
	reg  signed [ 9:0] r_sub05_V_addr;
	wire        [31:0] w_sub05_V_datain;
	reg         [31:0] r_sub05_V_datain;
	wire        [31:0] w_sub05_V_dataout;
	wire               w_sub05_V_r_w;
	reg                r_sub05_V_r_w;
	wire signed [ 9:0] w_sub05_U_addr;
	reg  signed [ 9:0] r_sub05_U_addr;
	wire        [31:0] w_sub05_U_datain;
	reg         [31:0] r_sub05_U_datain;
	wire        [31:0] w_sub05_U_dataout;
	wire               w_sub05_U_r_w;
	reg                r_sub05_U_r_w;
	wire signed [ 9:0] w_sub05_result_addr;
	reg  signed [ 9:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub18_run_req;
	wire               w_sub18_run_busy;
	wire signed [ 9:0] w_sub18_T_addr;
	reg  signed [ 9:0] r_sub18_T_addr;
	wire        [31:0] w_sub18_T_datain;
	reg         [31:0] r_sub18_T_datain;
	wire        [31:0] w_sub18_T_dataout;
	wire               w_sub18_T_r_w;
	reg                r_sub18_T_r_w;
	wire signed [ 9:0] w_sub18_V_addr;
	reg  signed [ 9:0] r_sub18_V_addr;
	wire        [31:0] w_sub18_V_datain;
	reg         [31:0] r_sub18_V_datain;
	wire        [31:0] w_sub18_V_dataout;
	wire               w_sub18_V_r_w;
	reg                r_sub18_V_r_w;
	wire signed [ 9:0] w_sub18_U_addr;
	reg  signed [ 9:0] r_sub18_U_addr;
	wire        [31:0] w_sub18_U_datain;
	reg         [31:0] r_sub18_U_datain;
	wire        [31:0] w_sub18_U_dataout;
	wire               w_sub18_U_r_w;
	reg                r_sub18_U_r_w;
	wire signed [ 9:0] w_sub18_result_addr;
	reg  signed [ 9:0] r_sub18_result_addr;
	wire        [31:0] w_sub18_result_datain;
	reg         [31:0] r_sub18_result_datain;
	wire        [31:0] w_sub18_result_dataout;
	wire               w_sub18_result_r_w;
	reg                r_sub18_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [ 9:0] w_sub04_T_addr;
	reg  signed [ 9:0] r_sub04_T_addr;
	wire        [31:0] w_sub04_T_datain;
	reg         [31:0] r_sub04_T_datain;
	wire        [31:0] w_sub04_T_dataout;
	wire               w_sub04_T_r_w;
	reg                r_sub04_T_r_w;
	wire signed [ 9:0] w_sub04_V_addr;
	reg  signed [ 9:0] r_sub04_V_addr;
	wire        [31:0] w_sub04_V_datain;
	reg         [31:0] r_sub04_V_datain;
	wire        [31:0] w_sub04_V_dataout;
	wire               w_sub04_V_r_w;
	reg                r_sub04_V_r_w;
	wire signed [ 9:0] w_sub04_U_addr;
	reg  signed [ 9:0] r_sub04_U_addr;
	wire        [31:0] w_sub04_U_datain;
	reg         [31:0] r_sub04_U_datain;
	wire        [31:0] w_sub04_U_dataout;
	wire               w_sub04_U_r_w;
	reg                r_sub04_U_r_w;
	wire signed [ 9:0] w_sub04_result_addr;
	reg  signed [ 9:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub17_run_req;
	wire               w_sub17_run_busy;
	wire signed [ 9:0] w_sub17_T_addr;
	reg  signed [ 9:0] r_sub17_T_addr;
	wire        [31:0] w_sub17_T_datain;
	reg         [31:0] r_sub17_T_datain;
	wire        [31:0] w_sub17_T_dataout;
	wire               w_sub17_T_r_w;
	reg                r_sub17_T_r_w;
	wire signed [ 9:0] w_sub17_V_addr;
	reg  signed [ 9:0] r_sub17_V_addr;
	wire        [31:0] w_sub17_V_datain;
	reg         [31:0] r_sub17_V_datain;
	wire        [31:0] w_sub17_V_dataout;
	wire               w_sub17_V_r_w;
	reg                r_sub17_V_r_w;
	wire signed [ 9:0] w_sub17_U_addr;
	reg  signed [ 9:0] r_sub17_U_addr;
	wire        [31:0] w_sub17_U_datain;
	reg         [31:0] r_sub17_U_datain;
	wire        [31:0] w_sub17_U_dataout;
	wire               w_sub17_U_r_w;
	reg                r_sub17_U_r_w;
	wire signed [ 9:0] w_sub17_result_addr;
	reg  signed [ 9:0] r_sub17_result_addr;
	wire        [31:0] w_sub17_result_datain;
	reg         [31:0] r_sub17_result_datain;
	wire        [31:0] w_sub17_result_dataout;
	wire               w_sub17_result_r_w;
	reg                r_sub17_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [ 9:0] w_sub10_T_addr;
	reg  signed [ 9:0] r_sub10_T_addr;
	wire        [31:0] w_sub10_T_datain;
	reg         [31:0] r_sub10_T_datain;
	wire        [31:0] w_sub10_T_dataout;
	wire               w_sub10_T_r_w;
	reg                r_sub10_T_r_w;
	wire signed [ 9:0] w_sub10_V_addr;
	reg  signed [ 9:0] r_sub10_V_addr;
	wire        [31:0] w_sub10_V_datain;
	reg         [31:0] r_sub10_V_datain;
	wire        [31:0] w_sub10_V_dataout;
	wire               w_sub10_V_r_w;
	reg                r_sub10_V_r_w;
	wire signed [ 9:0] w_sub10_U_addr;
	reg  signed [ 9:0] r_sub10_U_addr;
	wire        [31:0] w_sub10_U_datain;
	reg         [31:0] r_sub10_U_datain;
	wire        [31:0] w_sub10_U_dataout;
	wire               w_sub10_U_r_w;
	reg                r_sub10_U_r_w;
	wire signed [ 9:0] w_sub10_result_addr;
	reg  signed [ 9:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg                r_sub20_run_req;
	wire               w_sub20_run_busy;
	wire signed [ 9:0] w_sub20_T_addr;
	reg  signed [ 9:0] r_sub20_T_addr;
	wire        [31:0] w_sub20_T_datain;
	reg         [31:0] r_sub20_T_datain;
	wire        [31:0] w_sub20_T_dataout;
	wire               w_sub20_T_r_w;
	reg                r_sub20_T_r_w;
	wire signed [ 9:0] w_sub20_V_addr;
	reg  signed [ 9:0] r_sub20_V_addr;
	wire        [31:0] w_sub20_V_datain;
	reg         [31:0] r_sub20_V_datain;
	wire        [31:0] w_sub20_V_dataout;
	wire               w_sub20_V_r_w;
	reg                r_sub20_V_r_w;
	wire signed [ 9:0] w_sub20_U_addr;
	reg  signed [ 9:0] r_sub20_U_addr;
	wire        [31:0] w_sub20_U_datain;
	reg         [31:0] r_sub20_U_datain;
	wire        [31:0] w_sub20_U_dataout;
	wire               w_sub20_U_r_w;
	reg                r_sub20_U_r_w;
	wire signed [ 9:0] w_sub20_result_addr;
	reg  signed [ 9:0] r_sub20_result_addr;
	wire        [31:0] w_sub20_result_datain;
	reg         [31:0] r_sub20_result_datain;
	wire        [31:0] w_sub20_result_dataout;
	wire               w_sub20_result_r_w;
	reg                r_sub20_result_r_w;
	reg                r_sub21_run_req;
	wire               w_sub21_run_busy;
	wire signed [ 9:0] w_sub21_T_addr;
	reg  signed [ 9:0] r_sub21_T_addr;
	wire        [31:0] w_sub21_T_datain;
	reg         [31:0] r_sub21_T_datain;
	wire        [31:0] w_sub21_T_dataout;
	wire               w_sub21_T_r_w;
	reg                r_sub21_T_r_w;
	wire signed [ 9:0] w_sub21_V_addr;
	reg  signed [ 9:0] r_sub21_V_addr;
	wire        [31:0] w_sub21_V_datain;
	reg         [31:0] r_sub21_V_datain;
	wire        [31:0] w_sub21_V_dataout;
	wire               w_sub21_V_r_w;
	reg                r_sub21_V_r_w;
	wire signed [ 9:0] w_sub21_U_addr;
	reg  signed [ 9:0] r_sub21_U_addr;
	wire        [31:0] w_sub21_U_datain;
	reg         [31:0] r_sub21_U_datain;
	wire        [31:0] w_sub21_U_dataout;
	wire               w_sub21_U_r_w;
	reg                r_sub21_U_r_w;
	wire signed [ 9:0] w_sub21_result_addr;
	reg  signed [ 9:0] r_sub21_result_addr;
	wire        [31:0] w_sub21_result_datain;
	reg         [31:0] r_sub21_result_datain;
	wire        [31:0] w_sub21_result_dataout;
	wire               w_sub21_result_r_w;
	reg                r_sub21_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	reg         [31:0] r_sys_tmp48_float;
	reg         [31:0] r_sys_tmp49_float;
	reg         [31:0] r_sys_tmp50_float;
	reg         [31:0] r_sys_tmp51_float;
	reg         [31:0] r_sys_tmp52_float;
	reg         [31:0] r_sys_tmp53_float;
	reg         [31:0] r_sys_tmp54_float;
	reg         [31:0] r_sys_tmp55_float;
	reg         [31:0] r_sys_tmp56_float;
	reg         [31:0] r_sys_tmp57_float;
	reg         [31:0] r_sys_tmp58_float;
	reg         [31:0] r_sys_tmp59_float;
	reg         [31:0] r_sys_tmp60_float;
	reg         [31:0] r_sys_tmp61_float;
	reg         [31:0] r_sys_tmp62_float;
	reg         [31:0] r_sys_tmp63_float;
	reg         [31:0] r_sys_tmp64_float;
	reg         [31:0] r_sys_tmp65_float;
	reg         [31:0] r_sys_tmp66_float;
	reg         [31:0] r_sys_tmp67_float;
	reg         [31:0] r_sys_tmp68_float;
	reg         [31:0] r_sys_tmp69_float;
	reg         [31:0] r_sys_tmp70_float;
	reg         [31:0] r_sys_tmp71_float;
	reg         [31:0] r_sys_tmp72_float;
	reg         [31:0] r_sys_tmp73_float;
	reg         [31:0] r_sys_tmp74_float;
	reg         [31:0] r_sys_tmp75_float;
	reg         [31:0] r_sys_tmp76_float;
	reg         [31:0] r_sys_tmp77_float;
	reg         [31:0] r_sys_tmp78_float;
	reg         [31:0] r_sys_tmp79_float;
	reg         [31:0] r_sys_tmp80_float;
	reg         [31:0] r_sys_tmp81_float;
	reg         [31:0] r_sys_tmp82_float;
	reg         [31:0] r_sys_tmp83_float;
	reg         [31:0] r_sys_tmp84_float;
	reg         [31:0] r_sys_tmp85_float;
	reg         [31:0] r_sys_tmp86_float;
	reg         [31:0] r_sys_tmp87_float;
	reg         [31:0] r_sys_tmp88_float;
	reg         [31:0] r_sys_tmp89_float;
	reg         [31:0] r_sys_tmp90_float;
	reg         [31:0] r_sys_tmp91_float;
	reg         [31:0] r_sys_tmp92_float;
	reg         [31:0] r_sys_tmp93_float;
	reg         [31:0] r_sys_tmp94_float;
	reg         [31:0] r_sys_tmp95_float;
	reg         [31:0] r_sys_tmp96_float;
	reg         [31:0] r_sys_tmp97_float;
	reg         [31:0] r_sys_tmp98_float;
	reg         [31:0] r_sys_tmp99_float;
	reg         [31:0] r_sys_tmp100_float;
	reg         [31:0] r_sys_tmp101_float;
	reg         [31:0] r_sys_tmp102_float;
	reg         [31:0] r_sys_tmp103_float;
	reg         [31:0] r_sys_tmp104_float;
	reg         [31:0] r_sys_tmp105_float;
	reg         [31:0] r_sys_tmp106_float;
	reg         [31:0] r_sys_tmp107_float;
	reg         [31:0] r_sys_tmp108_float;
	reg         [31:0] r_sys_tmp109_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire               w_sys_tmp12;
	wire               w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp15;
	wire               w_sys_tmp16;
	wire        [31:0] w_sys_tmp18;
	wire        [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire        [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp27;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp32;
	wire signed [31:0] w_sys_tmp33;
	wire        [31:0] w_sys_tmp36;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp45;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire        [31:0] w_sys_tmp128;
	wire               w_sys_tmp226;
	wire               w_sys_tmp227;
	wire signed [31:0] w_sys_tmp228;
	wire signed [31:0] w_sys_tmp231;
	wire signed [31:0] w_sys_tmp232;
	wire        [31:0] w_sys_tmp233;
	wire        [31:0] w_sys_tmp239;
	wire signed [31:0] w_sys_tmp243;
	wire signed [31:0] w_sys_tmp244;
	wire signed [31:0] w_sys_tmp255;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp267;
	wire signed [31:0] w_sys_tmp268;
	wire signed [31:0] w_sys_tmp279;
	wire signed [31:0] w_sys_tmp280;
	wire signed [31:0] w_sys_tmp291;
	wire signed [31:0] w_sys_tmp292;
	wire signed [31:0] w_sys_tmp303;
	wire signed [31:0] w_sys_tmp304;
	wire signed [31:0] w_sys_tmp315;
	wire signed [31:0] w_sys_tmp316;
	wire signed [31:0] w_sys_tmp351;
	wire signed [31:0] w_sys_tmp352;
	wire signed [31:0] w_sys_tmp363;
	wire signed [31:0] w_sys_tmp364;
	wire signed [31:0] w_sys_tmp375;
	wire signed [31:0] w_sys_tmp376;
	wire signed [31:0] w_sys_tmp387;
	wire signed [31:0] w_sys_tmp388;
	wire signed [31:0] w_sys_tmp399;
	wire signed [31:0] w_sys_tmp400;
	wire signed [31:0] w_sys_tmp411;
	wire signed [31:0] w_sys_tmp412;
	wire signed [31:0] w_sys_tmp447;
	wire signed [31:0] w_sys_tmp448;
	wire signed [31:0] w_sys_tmp459;
	wire signed [31:0] w_sys_tmp460;
	wire signed [31:0] w_sys_tmp471;
	wire signed [31:0] w_sys_tmp472;
	wire signed [31:0] w_sys_tmp483;
	wire signed [31:0] w_sys_tmp484;
	wire signed [31:0] w_sys_tmp495;
	wire signed [31:0] w_sys_tmp496;
	wire signed [31:0] w_sys_tmp507;
	wire signed [31:0] w_sys_tmp508;
	wire signed [31:0] w_sys_tmp543;
	wire signed [31:0] w_sys_tmp544;
	wire signed [31:0] w_sys_tmp555;
	wire signed [31:0] w_sys_tmp556;
	wire signed [31:0] w_sys_tmp567;
	wire signed [31:0] w_sys_tmp568;
	wire signed [31:0] w_sys_tmp579;
	wire signed [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp591;
	wire signed [31:0] w_sys_tmp592;
	wire signed [31:0] w_sys_tmp603;
	wire signed [31:0] w_sys_tmp604;
	wire signed [31:0] w_sys_tmp639;
	wire signed [31:0] w_sys_tmp640;
	wire signed [31:0] w_sys_tmp651;
	wire signed [31:0] w_sys_tmp652;
	wire signed [31:0] w_sys_tmp663;
	wire signed [31:0] w_sys_tmp664;
	wire signed [31:0] w_sys_tmp675;
	wire signed [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp687;
	wire signed [31:0] w_sys_tmp688;
	wire signed [31:0] w_sys_tmp699;
	wire signed [31:0] w_sys_tmp700;
	wire signed [31:0] w_sys_tmp711;
	wire signed [31:0] w_sys_tmp712;
	wire signed [31:0] w_sys_tmp723;
	wire signed [31:0] w_sys_tmp724;
	wire signed [31:0] w_sys_tmp735;
	wire signed [31:0] w_sys_tmp736;
	wire signed [31:0] w_sys_tmp747;
	wire signed [31:0] w_sys_tmp748;
	wire signed [31:0] w_sys_tmp759;
	wire signed [31:0] w_sys_tmp760;
	wire signed [31:0] w_sys_tmp771;
	wire signed [31:0] w_sys_tmp772;
	wire signed [31:0] w_sys_tmp783;
	wire signed [31:0] w_sys_tmp784;
	wire signed [31:0] w_sys_tmp819;
	wire signed [31:0] w_sys_tmp820;
	wire signed [31:0] w_sys_tmp831;
	wire signed [31:0] w_sys_tmp832;
	wire signed [31:0] w_sys_tmp843;
	wire signed [31:0] w_sys_tmp844;
	wire signed [31:0] w_sys_tmp855;
	wire signed [31:0] w_sys_tmp856;
	wire signed [31:0] w_sys_tmp867;
	wire signed [31:0] w_sys_tmp868;
	wire signed [31:0] w_sys_tmp879;
	wire signed [31:0] w_sys_tmp880;
	wire signed [31:0] w_sys_tmp915;
	wire signed [31:0] w_sys_tmp916;
	wire signed [31:0] w_sys_tmp927;
	wire signed [31:0] w_sys_tmp928;
	wire signed [31:0] w_sys_tmp939;
	wire signed [31:0] w_sys_tmp940;
	wire signed [31:0] w_sys_tmp951;
	wire signed [31:0] w_sys_tmp952;
	wire signed [31:0] w_sys_tmp963;
	wire signed [31:0] w_sys_tmp964;
	wire signed [31:0] w_sys_tmp975;
	wire signed [31:0] w_sys_tmp976;
	wire signed [31:0] w_sys_tmp1011;
	wire signed [31:0] w_sys_tmp1012;
	wire signed [31:0] w_sys_tmp1023;
	wire signed [31:0] w_sys_tmp1024;
	wire signed [31:0] w_sys_tmp1035;
	wire signed [31:0] w_sys_tmp1036;
	wire signed [31:0] w_sys_tmp1047;
	wire signed [31:0] w_sys_tmp1048;
	wire signed [31:0] w_sys_tmp1059;
	wire signed [31:0] w_sys_tmp1060;
	wire signed [31:0] w_sys_tmp1071;
	wire signed [31:0] w_sys_tmp1072;
	wire signed [31:0] w_sys_tmp1107;
	wire signed [31:0] w_sys_tmp1108;
	wire signed [31:0] w_sys_tmp1119;
	wire signed [31:0] w_sys_tmp1120;
	wire signed [31:0] w_sys_tmp1131;
	wire signed [31:0] w_sys_tmp1132;
	wire signed [31:0] w_sys_tmp1143;
	wire signed [31:0] w_sys_tmp1144;
	wire signed [31:0] w_sys_tmp1155;
	wire signed [31:0] w_sys_tmp1156;
	wire signed [31:0] w_sys_tmp1167;
	wire signed [31:0] w_sys_tmp1168;
	wire signed [31:0] w_sys_tmp1179;
	wire signed [31:0] w_sys_tmp1180;
	wire signed [31:0] w_sys_tmp1191;
	wire signed [31:0] w_sys_tmp1192;
	wire signed [31:0] w_sys_tmp1203;
	wire signed [31:0] w_sys_tmp1204;
	wire signed [31:0] w_sys_tmp1215;
	wire signed [31:0] w_sys_tmp1216;
	wire signed [31:0] w_sys_tmp1227;
	wire signed [31:0] w_sys_tmp1228;
	wire signed [31:0] w_sys_tmp1239;
	wire signed [31:0] w_sys_tmp1240;
	wire signed [31:0] w_sys_tmp1251;
	wire signed [31:0] w_sys_tmp1252;
	wire signed [31:0] w_sys_tmp1287;
	wire signed [31:0] w_sys_tmp1288;
	wire signed [31:0] w_sys_tmp1299;
	wire signed [31:0] w_sys_tmp1300;
	wire signed [31:0] w_sys_tmp1311;
	wire signed [31:0] w_sys_tmp1312;
	wire signed [31:0] w_sys_tmp1323;
	wire signed [31:0] w_sys_tmp1324;
	wire signed [31:0] w_sys_tmp1335;
	wire signed [31:0] w_sys_tmp1336;
	wire signed [31:0] w_sys_tmp1347;
	wire signed [31:0] w_sys_tmp1348;
	wire signed [31:0] w_sys_tmp1383;
	wire signed [31:0] w_sys_tmp1384;
	wire signed [31:0] w_sys_tmp1395;
	wire signed [31:0] w_sys_tmp1396;
	wire signed [31:0] w_sys_tmp1407;
	wire signed [31:0] w_sys_tmp1408;
	wire signed [31:0] w_sys_tmp1419;
	wire signed [31:0] w_sys_tmp1420;
	wire signed [31:0] w_sys_tmp1431;
	wire signed [31:0] w_sys_tmp1432;
	wire signed [31:0] w_sys_tmp1443;
	wire signed [31:0] w_sys_tmp1444;
	wire signed [31:0] w_sys_tmp1479;
	wire signed [31:0] w_sys_tmp1480;
	wire signed [31:0] w_sys_tmp1491;
	wire signed [31:0] w_sys_tmp1492;
	wire signed [31:0] w_sys_tmp1503;
	wire signed [31:0] w_sys_tmp1504;
	wire signed [31:0] w_sys_tmp1515;
	wire signed [31:0] w_sys_tmp1516;
	wire signed [31:0] w_sys_tmp1527;
	wire signed [31:0] w_sys_tmp1528;
	wire signed [31:0] w_sys_tmp1539;
	wire signed [31:0] w_sys_tmp1540;
	wire signed [31:0] w_sys_tmp1575;
	wire signed [31:0] w_sys_tmp1576;
	wire signed [31:0] w_sys_tmp1587;
	wire signed [31:0] w_sys_tmp1588;
	wire signed [31:0] w_sys_tmp1599;
	wire signed [31:0] w_sys_tmp1600;
	wire signed [31:0] w_sys_tmp1611;
	wire signed [31:0] w_sys_tmp1612;
	wire signed [31:0] w_sys_tmp1623;
	wire signed [31:0] w_sys_tmp1624;
	wire signed [31:0] w_sys_tmp1635;
	wire signed [31:0] w_sys_tmp1636;
	wire signed [31:0] w_sys_tmp1647;
	wire signed [31:0] w_sys_tmp1648;
	wire signed [31:0] w_sys_tmp1659;
	wire signed [31:0] w_sys_tmp1660;
	wire signed [31:0] w_sys_tmp1671;
	wire signed [31:0] w_sys_tmp1672;
	wire signed [31:0] w_sys_tmp1683;
	wire signed [31:0] w_sys_tmp1684;
	wire signed [31:0] w_sys_tmp1695;
	wire signed [31:0] w_sys_tmp1696;
	wire signed [31:0] w_sys_tmp1707;
	wire signed [31:0] w_sys_tmp1708;
	wire signed [31:0] w_sys_tmp1719;
	wire signed [31:0] w_sys_tmp1720;
	wire signed [31:0] w_sys_tmp1755;
	wire signed [31:0] w_sys_tmp1756;
	wire signed [31:0] w_sys_tmp1767;
	wire signed [31:0] w_sys_tmp1768;
	wire signed [31:0] w_sys_tmp1779;
	wire signed [31:0] w_sys_tmp1780;
	wire signed [31:0] w_sys_tmp1791;
	wire signed [31:0] w_sys_tmp1792;
	wire signed [31:0] w_sys_tmp1803;
	wire signed [31:0] w_sys_tmp1804;
	wire signed [31:0] w_sys_tmp1815;
	wire signed [31:0] w_sys_tmp1816;
	wire signed [31:0] w_sys_tmp1851;
	wire signed [31:0] w_sys_tmp1852;
	wire signed [31:0] w_sys_tmp1863;
	wire signed [31:0] w_sys_tmp1864;
	wire signed [31:0] w_sys_tmp1875;
	wire signed [31:0] w_sys_tmp1876;
	wire signed [31:0] w_sys_tmp1887;
	wire signed [31:0] w_sys_tmp1888;
	wire signed [31:0] w_sys_tmp1899;
	wire signed [31:0] w_sys_tmp1900;
	wire signed [31:0] w_sys_tmp1911;
	wire signed [31:0] w_sys_tmp1912;
	wire signed [31:0] w_sys_tmp1947;
	wire signed [31:0] w_sys_tmp1948;
	wire signed [31:0] w_sys_tmp1959;
	wire signed [31:0] w_sys_tmp1960;
	wire signed [31:0] w_sys_tmp1971;
	wire signed [31:0] w_sys_tmp1972;
	wire signed [31:0] w_sys_tmp1983;
	wire signed [31:0] w_sys_tmp1984;
	wire signed [31:0] w_sys_tmp1995;
	wire signed [31:0] w_sys_tmp1996;
	wire signed [31:0] w_sys_tmp2007;
	wire signed [31:0] w_sys_tmp2008;
	wire signed [31:0] w_sys_tmp2043;
	wire signed [31:0] w_sys_tmp2044;
	wire signed [31:0] w_sys_tmp2055;
	wire signed [31:0] w_sys_tmp2056;
	wire signed [31:0] w_sys_tmp2067;
	wire signed [31:0] w_sys_tmp2068;
	wire signed [31:0] w_sys_tmp2079;
	wire signed [31:0] w_sys_tmp2080;
	wire signed [31:0] w_sys_tmp2091;
	wire signed [31:0] w_sys_tmp2092;
	wire signed [31:0] w_sys_tmp2102;
	wire signed [31:0] w_sys_tmp2103;
	wire               w_sys_tmp2104;
	wire               w_sys_tmp2105;
	wire signed [31:0] w_sys_tmp2106;
	wire signed [31:0] w_sys_tmp2109;
	wire signed [31:0] w_sys_tmp2110;
	wire        [31:0] w_sys_tmp2111;
	wire        [31:0] w_sys_tmp2117;
	wire signed [31:0] w_sys_tmp2121;
	wire signed [31:0] w_sys_tmp2122;
	wire signed [31:0] w_sys_tmp2133;
	wire signed [31:0] w_sys_tmp2134;
	wire signed [31:0] w_sys_tmp2145;
	wire signed [31:0] w_sys_tmp2146;
	wire signed [31:0] w_sys_tmp2157;
	wire signed [31:0] w_sys_tmp2158;
	wire signed [31:0] w_sys_tmp2169;
	wire signed [31:0] w_sys_tmp2170;
	wire signed [31:0] w_sys_tmp2181;
	wire signed [31:0] w_sys_tmp2182;
	wire signed [31:0] w_sys_tmp2193;
	wire signed [31:0] w_sys_tmp2194;
	wire signed [31:0] w_sys_tmp2229;
	wire signed [31:0] w_sys_tmp2230;
	wire signed [31:0] w_sys_tmp2241;
	wire signed [31:0] w_sys_tmp2242;
	wire signed [31:0] w_sys_tmp2253;
	wire signed [31:0] w_sys_tmp2254;
	wire signed [31:0] w_sys_tmp2265;
	wire signed [31:0] w_sys_tmp2266;
	wire signed [31:0] w_sys_tmp2277;
	wire signed [31:0] w_sys_tmp2278;
	wire signed [31:0] w_sys_tmp2289;
	wire signed [31:0] w_sys_tmp2290;
	wire signed [31:0] w_sys_tmp2325;
	wire signed [31:0] w_sys_tmp2326;
	wire signed [31:0] w_sys_tmp2337;
	wire signed [31:0] w_sys_tmp2338;
	wire signed [31:0] w_sys_tmp2349;
	wire signed [31:0] w_sys_tmp2350;
	wire signed [31:0] w_sys_tmp2361;
	wire signed [31:0] w_sys_tmp2362;
	wire signed [31:0] w_sys_tmp2373;
	wire signed [31:0] w_sys_tmp2374;
	wire signed [31:0] w_sys_tmp2385;
	wire signed [31:0] w_sys_tmp2386;
	wire signed [31:0] w_sys_tmp2421;
	wire signed [31:0] w_sys_tmp2422;
	wire signed [31:0] w_sys_tmp2433;
	wire signed [31:0] w_sys_tmp2434;
	wire signed [31:0] w_sys_tmp2445;
	wire signed [31:0] w_sys_tmp2446;
	wire signed [31:0] w_sys_tmp2457;
	wire signed [31:0] w_sys_tmp2458;
	wire signed [31:0] w_sys_tmp2469;
	wire signed [31:0] w_sys_tmp2470;
	wire signed [31:0] w_sys_tmp2481;
	wire signed [31:0] w_sys_tmp2482;
	wire signed [31:0] w_sys_tmp2517;
	wire signed [31:0] w_sys_tmp2518;
	wire signed [31:0] w_sys_tmp2529;
	wire signed [31:0] w_sys_tmp2530;
	wire signed [31:0] w_sys_tmp2541;
	wire signed [31:0] w_sys_tmp2542;
	wire signed [31:0] w_sys_tmp2553;
	wire signed [31:0] w_sys_tmp2554;
	wire signed [31:0] w_sys_tmp2565;
	wire signed [31:0] w_sys_tmp2566;
	wire signed [31:0] w_sys_tmp2576;
	wire               w_sys_tmp2577;
	wire               w_sys_tmp2578;
	wire signed [31:0] w_sys_tmp2579;
	wire               w_sys_tmp2580;
	wire               w_sys_tmp2581;
	wire signed [31:0] w_sys_tmp2584;
	wire signed [31:0] w_sys_tmp2585;
	wire        [31:0] w_sys_tmp2586;
	wire signed [31:0] w_sys_tmp2588;
	wire signed [31:0] w_sys_tmp2589;
	wire        [31:0] w_sys_tmp2591;
	wire signed [31:0] w_sys_tmp2592;
	wire signed [31:0] w_sys_tmp2593;
	wire signed [31:0] w_sys_tmp2594;
	wire signed [31:0] w_sys_tmp2596;
	wire               w_sys_tmp2597;
	wire               w_sys_tmp2598;
	wire signed [31:0] w_sys_tmp2601;
	wire signed [31:0] w_sys_tmp2602;
	wire signed [31:0] w_sys_tmp2603;
	wire        [31:0] w_sys_tmp2604;
	wire signed [31:0] w_sys_tmp2606;
	wire signed [31:0] w_sys_tmp2607;
	wire signed [31:0] w_sys_tmp2610;
	wire signed [31:0] w_sys_tmp2611;
	wire signed [31:0] w_sys_tmp2684;
	wire signed [31:0] w_sys_tmp2685;
	wire               w_sys_tmp2686;
	wire               w_sys_tmp2687;
	wire signed [31:0] w_sys_tmp2688;
	wire signed [31:0] w_sys_tmp2689;
	wire signed [31:0] w_sys_tmp2692;
	wire signed [31:0] w_sys_tmp2693;
	wire signed [31:0] w_sys_tmp2694;
	wire        [31:0] w_sys_tmp2695;
	wire signed [31:0] w_sys_tmp2696;
	wire               w_sys_tmp2733;
	wire               w_sys_tmp2734;
	wire signed [31:0] w_sys_tmp2735;
	wire signed [31:0] w_sys_tmp2738;
	wire signed [31:0] w_sys_tmp2739;
	wire        [31:0] w_sys_tmp2740;
	wire signed [31:0] w_sys_tmp2744;
	wire signed [31:0] w_sys_tmp2745;
	wire signed [31:0] w_sys_tmp2750;
	wire signed [31:0] w_sys_tmp2751;
	wire signed [31:0] w_sys_tmp2756;
	wire signed [31:0] w_sys_tmp2757;
	wire signed [31:0] w_sys_tmp2762;
	wire signed [31:0] w_sys_tmp2763;
	wire signed [31:0] w_sys_tmp2768;
	wire signed [31:0] w_sys_tmp2769;
	wire signed [31:0] w_sys_tmp2774;
	wire signed [31:0] w_sys_tmp2775;
	wire signed [31:0] w_sys_tmp2780;
	wire signed [31:0] w_sys_tmp2781;
	wire signed [31:0] w_sys_tmp2798;
	wire signed [31:0] w_sys_tmp2799;
	wire signed [31:0] w_sys_tmp2804;
	wire signed [31:0] w_sys_tmp2805;
	wire signed [31:0] w_sys_tmp2810;
	wire signed [31:0] w_sys_tmp2811;
	wire signed [31:0] w_sys_tmp2816;
	wire signed [31:0] w_sys_tmp2817;
	wire signed [31:0] w_sys_tmp2822;
	wire signed [31:0] w_sys_tmp2823;
	wire signed [31:0] w_sys_tmp2828;
	wire signed [31:0] w_sys_tmp2829;
	wire signed [31:0] w_sys_tmp2846;
	wire signed [31:0] w_sys_tmp2847;
	wire signed [31:0] w_sys_tmp2852;
	wire signed [31:0] w_sys_tmp2853;
	wire signed [31:0] w_sys_tmp2858;
	wire signed [31:0] w_sys_tmp2859;
	wire signed [31:0] w_sys_tmp2864;
	wire signed [31:0] w_sys_tmp2865;
	wire signed [31:0] w_sys_tmp2870;
	wire signed [31:0] w_sys_tmp2871;
	wire signed [31:0] w_sys_tmp2876;
	wire signed [31:0] w_sys_tmp2877;
	wire signed [31:0] w_sys_tmp2894;
	wire signed [31:0] w_sys_tmp2895;
	wire signed [31:0] w_sys_tmp2900;
	wire signed [31:0] w_sys_tmp2901;
	wire signed [31:0] w_sys_tmp2906;
	wire signed [31:0] w_sys_tmp2907;
	wire signed [31:0] w_sys_tmp2912;
	wire signed [31:0] w_sys_tmp2913;
	wire signed [31:0] w_sys_tmp2918;
	wire signed [31:0] w_sys_tmp2919;
	wire signed [31:0] w_sys_tmp2924;
	wire signed [31:0] w_sys_tmp2925;
	wire signed [31:0] w_sys_tmp2942;
	wire signed [31:0] w_sys_tmp2943;
	wire signed [31:0] w_sys_tmp2948;
	wire signed [31:0] w_sys_tmp2949;
	wire signed [31:0] w_sys_tmp2954;
	wire signed [31:0] w_sys_tmp2955;
	wire signed [31:0] w_sys_tmp2960;
	wire signed [31:0] w_sys_tmp2961;
	wire signed [31:0] w_sys_tmp2966;
	wire signed [31:0] w_sys_tmp2967;
	wire signed [31:0] w_sys_tmp2972;
	wire signed [31:0] w_sys_tmp2973;
	wire signed [31:0] w_sys_tmp2978;
	wire signed [31:0] w_sys_tmp2979;
	wire signed [31:0] w_sys_tmp2984;
	wire signed [31:0] w_sys_tmp2985;
	wire signed [31:0] w_sys_tmp2990;
	wire signed [31:0] w_sys_tmp2991;
	wire signed [31:0] w_sys_tmp2996;
	wire signed [31:0] w_sys_tmp2997;
	wire signed [31:0] w_sys_tmp3002;
	wire signed [31:0] w_sys_tmp3003;
	wire signed [31:0] w_sys_tmp3008;
	wire signed [31:0] w_sys_tmp3009;
	wire signed [31:0] w_sys_tmp3014;
	wire signed [31:0] w_sys_tmp3015;
	wire signed [31:0] w_sys_tmp3032;
	wire signed [31:0] w_sys_tmp3033;
	wire signed [31:0] w_sys_tmp3038;
	wire signed [31:0] w_sys_tmp3039;
	wire signed [31:0] w_sys_tmp3044;
	wire signed [31:0] w_sys_tmp3045;
	wire signed [31:0] w_sys_tmp3050;
	wire signed [31:0] w_sys_tmp3051;
	wire signed [31:0] w_sys_tmp3056;
	wire signed [31:0] w_sys_tmp3057;
	wire signed [31:0] w_sys_tmp3062;
	wire signed [31:0] w_sys_tmp3063;
	wire signed [31:0] w_sys_tmp3080;
	wire signed [31:0] w_sys_tmp3081;
	wire signed [31:0] w_sys_tmp3086;
	wire signed [31:0] w_sys_tmp3087;
	wire signed [31:0] w_sys_tmp3092;
	wire signed [31:0] w_sys_tmp3093;
	wire signed [31:0] w_sys_tmp3098;
	wire signed [31:0] w_sys_tmp3099;
	wire signed [31:0] w_sys_tmp3104;
	wire signed [31:0] w_sys_tmp3105;
	wire signed [31:0] w_sys_tmp3110;
	wire signed [31:0] w_sys_tmp3111;
	wire signed [31:0] w_sys_tmp3128;
	wire signed [31:0] w_sys_tmp3129;
	wire signed [31:0] w_sys_tmp3134;
	wire signed [31:0] w_sys_tmp3135;
	wire signed [31:0] w_sys_tmp3140;
	wire signed [31:0] w_sys_tmp3141;
	wire signed [31:0] w_sys_tmp3146;
	wire signed [31:0] w_sys_tmp3147;
	wire signed [31:0] w_sys_tmp3152;
	wire signed [31:0] w_sys_tmp3153;
	wire signed [31:0] w_sys_tmp3158;
	wire signed [31:0] w_sys_tmp3159;
	wire signed [31:0] w_sys_tmp3176;
	wire signed [31:0] w_sys_tmp3177;
	wire signed [31:0] w_sys_tmp3182;
	wire signed [31:0] w_sys_tmp3183;
	wire signed [31:0] w_sys_tmp3188;
	wire signed [31:0] w_sys_tmp3189;
	wire signed [31:0] w_sys_tmp3194;
	wire signed [31:0] w_sys_tmp3195;
	wire signed [31:0] w_sys_tmp3200;
	wire signed [31:0] w_sys_tmp3201;
	wire signed [31:0] w_sys_tmp3206;
	wire signed [31:0] w_sys_tmp3207;
	wire signed [31:0] w_sys_tmp3212;
	wire signed [31:0] w_sys_tmp3213;
	wire signed [31:0] w_sys_tmp3218;
	wire signed [31:0] w_sys_tmp3219;
	wire signed [31:0] w_sys_tmp3224;
	wire signed [31:0] w_sys_tmp3225;
	wire signed [31:0] w_sys_tmp3230;
	wire signed [31:0] w_sys_tmp3231;
	wire signed [31:0] w_sys_tmp3236;
	wire signed [31:0] w_sys_tmp3237;
	wire signed [31:0] w_sys_tmp3242;
	wire signed [31:0] w_sys_tmp3243;
	wire signed [31:0] w_sys_tmp3248;
	wire signed [31:0] w_sys_tmp3249;
	wire signed [31:0] w_sys_tmp3266;
	wire signed [31:0] w_sys_tmp3267;
	wire signed [31:0] w_sys_tmp3272;
	wire signed [31:0] w_sys_tmp3273;
	wire signed [31:0] w_sys_tmp3278;
	wire signed [31:0] w_sys_tmp3279;
	wire signed [31:0] w_sys_tmp3284;
	wire signed [31:0] w_sys_tmp3285;
	wire signed [31:0] w_sys_tmp3290;
	wire signed [31:0] w_sys_tmp3291;
	wire signed [31:0] w_sys_tmp3296;
	wire signed [31:0] w_sys_tmp3297;
	wire signed [31:0] w_sys_tmp3314;
	wire signed [31:0] w_sys_tmp3315;
	wire signed [31:0] w_sys_tmp3320;
	wire signed [31:0] w_sys_tmp3321;
	wire signed [31:0] w_sys_tmp3326;
	wire signed [31:0] w_sys_tmp3327;
	wire signed [31:0] w_sys_tmp3332;
	wire signed [31:0] w_sys_tmp3333;
	wire signed [31:0] w_sys_tmp3338;
	wire signed [31:0] w_sys_tmp3339;
	wire signed [31:0] w_sys_tmp3344;
	wire signed [31:0] w_sys_tmp3345;
	wire signed [31:0] w_sys_tmp3362;
	wire signed [31:0] w_sys_tmp3363;
	wire signed [31:0] w_sys_tmp3368;
	wire signed [31:0] w_sys_tmp3369;
	wire signed [31:0] w_sys_tmp3374;
	wire signed [31:0] w_sys_tmp3375;
	wire signed [31:0] w_sys_tmp3380;
	wire signed [31:0] w_sys_tmp3381;
	wire signed [31:0] w_sys_tmp3386;
	wire signed [31:0] w_sys_tmp3387;
	wire signed [31:0] w_sys_tmp3392;
	wire signed [31:0] w_sys_tmp3393;
	wire signed [31:0] w_sys_tmp3410;
	wire signed [31:0] w_sys_tmp3411;
	wire signed [31:0] w_sys_tmp3416;
	wire signed [31:0] w_sys_tmp3417;
	wire signed [31:0] w_sys_tmp3422;
	wire signed [31:0] w_sys_tmp3423;
	wire signed [31:0] w_sys_tmp3428;
	wire signed [31:0] w_sys_tmp3429;
	wire signed [31:0] w_sys_tmp3434;
	wire signed [31:0] w_sys_tmp3435;
	wire signed [31:0] w_sys_tmp3440;
	wire signed [31:0] w_sys_tmp3441;
	wire signed [31:0] w_sys_tmp3446;
	wire signed [31:0] w_sys_tmp3447;
	wire signed [31:0] w_sys_tmp3452;
	wire signed [31:0] w_sys_tmp3453;
	wire signed [31:0] w_sys_tmp3458;
	wire signed [31:0] w_sys_tmp3459;
	wire signed [31:0] w_sys_tmp3464;
	wire signed [31:0] w_sys_tmp3465;
	wire signed [31:0] w_sys_tmp3470;
	wire signed [31:0] w_sys_tmp3471;
	wire signed [31:0] w_sys_tmp3476;
	wire signed [31:0] w_sys_tmp3477;
	wire signed [31:0] w_sys_tmp3482;
	wire signed [31:0] w_sys_tmp3483;
	wire signed [31:0] w_sys_tmp3500;
	wire signed [31:0] w_sys_tmp3501;
	wire signed [31:0] w_sys_tmp3506;
	wire signed [31:0] w_sys_tmp3507;
	wire signed [31:0] w_sys_tmp3512;
	wire signed [31:0] w_sys_tmp3513;
	wire signed [31:0] w_sys_tmp3518;
	wire signed [31:0] w_sys_tmp3519;
	wire signed [31:0] w_sys_tmp3524;
	wire signed [31:0] w_sys_tmp3525;
	wire signed [31:0] w_sys_tmp3530;
	wire signed [31:0] w_sys_tmp3531;
	wire signed [31:0] w_sys_tmp3548;
	wire signed [31:0] w_sys_tmp3549;
	wire signed [31:0] w_sys_tmp3554;
	wire signed [31:0] w_sys_tmp3555;
	wire signed [31:0] w_sys_tmp3560;
	wire signed [31:0] w_sys_tmp3561;
	wire signed [31:0] w_sys_tmp3566;
	wire signed [31:0] w_sys_tmp3567;
	wire signed [31:0] w_sys_tmp3572;
	wire signed [31:0] w_sys_tmp3573;
	wire signed [31:0] w_sys_tmp3578;
	wire signed [31:0] w_sys_tmp3579;
	wire signed [31:0] w_sys_tmp3596;
	wire signed [31:0] w_sys_tmp3597;
	wire signed [31:0] w_sys_tmp3602;
	wire signed [31:0] w_sys_tmp3603;
	wire signed [31:0] w_sys_tmp3608;
	wire signed [31:0] w_sys_tmp3609;
	wire signed [31:0] w_sys_tmp3614;
	wire signed [31:0] w_sys_tmp3615;
	wire signed [31:0] w_sys_tmp3620;
	wire signed [31:0] w_sys_tmp3621;
	wire signed [31:0] w_sys_tmp3626;
	wire signed [31:0] w_sys_tmp3627;
	wire signed [31:0] w_sys_tmp3644;
	wire signed [31:0] w_sys_tmp3645;
	wire signed [31:0] w_sys_tmp3650;
	wire signed [31:0] w_sys_tmp3651;
	wire signed [31:0] w_sys_tmp3656;
	wire signed [31:0] w_sys_tmp3657;
	wire signed [31:0] w_sys_tmp3662;
	wire signed [31:0] w_sys_tmp3663;
	wire signed [31:0] w_sys_tmp3668;
	wire signed [31:0] w_sys_tmp3669;
	wire signed [31:0] w_sys_tmp3673;
	wire signed [31:0] w_sys_tmp3674;
	wire               w_sys_tmp3675;
	wire               w_sys_tmp3676;
	wire signed [31:0] w_sys_tmp3677;
	wire signed [31:0] w_sys_tmp3680;
	wire signed [31:0] w_sys_tmp3681;
	wire        [31:0] w_sys_tmp3682;
	wire signed [31:0] w_sys_tmp3686;
	wire signed [31:0] w_sys_tmp3687;
	wire signed [31:0] w_sys_tmp3692;
	wire signed [31:0] w_sys_tmp3693;
	wire signed [31:0] w_sys_tmp3698;
	wire signed [31:0] w_sys_tmp3699;
	wire signed [31:0] w_sys_tmp3704;
	wire signed [31:0] w_sys_tmp3705;
	wire signed [31:0] w_sys_tmp3710;
	wire signed [31:0] w_sys_tmp3711;
	wire signed [31:0] w_sys_tmp3716;
	wire signed [31:0] w_sys_tmp3717;
	wire signed [31:0] w_sys_tmp3722;
	wire signed [31:0] w_sys_tmp3723;
	wire signed [31:0] w_sys_tmp3740;
	wire signed [31:0] w_sys_tmp3741;
	wire signed [31:0] w_sys_tmp3746;
	wire signed [31:0] w_sys_tmp3747;
	wire signed [31:0] w_sys_tmp3752;
	wire signed [31:0] w_sys_tmp3753;
	wire signed [31:0] w_sys_tmp3758;
	wire signed [31:0] w_sys_tmp3759;
	wire signed [31:0] w_sys_tmp3764;
	wire signed [31:0] w_sys_tmp3765;
	wire signed [31:0] w_sys_tmp3770;
	wire signed [31:0] w_sys_tmp3771;
	wire signed [31:0] w_sys_tmp3788;
	wire signed [31:0] w_sys_tmp3789;
	wire signed [31:0] w_sys_tmp3794;
	wire signed [31:0] w_sys_tmp3795;
	wire signed [31:0] w_sys_tmp3800;
	wire signed [31:0] w_sys_tmp3801;
	wire signed [31:0] w_sys_tmp3806;
	wire signed [31:0] w_sys_tmp3807;
	wire signed [31:0] w_sys_tmp3812;
	wire signed [31:0] w_sys_tmp3813;
	wire signed [31:0] w_sys_tmp3818;
	wire signed [31:0] w_sys_tmp3819;
	wire signed [31:0] w_sys_tmp3836;
	wire signed [31:0] w_sys_tmp3837;
	wire signed [31:0] w_sys_tmp3842;
	wire signed [31:0] w_sys_tmp3843;
	wire signed [31:0] w_sys_tmp3848;
	wire signed [31:0] w_sys_tmp3849;
	wire signed [31:0] w_sys_tmp3854;
	wire signed [31:0] w_sys_tmp3855;
	wire signed [31:0] w_sys_tmp3860;
	wire signed [31:0] w_sys_tmp3861;
	wire signed [31:0] w_sys_tmp3866;
	wire signed [31:0] w_sys_tmp3867;
	wire signed [31:0] w_sys_tmp3884;
	wire signed [31:0] w_sys_tmp3885;
	wire signed [31:0] w_sys_tmp3890;
	wire signed [31:0] w_sys_tmp3891;
	wire signed [31:0] w_sys_tmp3896;
	wire signed [31:0] w_sys_tmp3897;
	wire signed [31:0] w_sys_tmp3902;
	wire signed [31:0] w_sys_tmp3903;
	wire signed [31:0] w_sys_tmp3908;
	wire signed [31:0] w_sys_tmp3909;
	wire signed [31:0] w_sys_tmp3913;
	wire signed [31:0] w_sys_tmp3914;
	wire               w_sys_tmp3915;
	wire               w_sys_tmp3916;
	wire signed [31:0] w_sys_tmp3917;
	wire signed [31:0] w_sys_tmp3920;
	wire signed [31:0] w_sys_tmp3921;
	wire        [31:0] w_sys_tmp3922;
	wire signed [31:0] w_sys_tmp3926;
	wire signed [31:0] w_sys_tmp3927;
	wire signed [31:0] w_sys_tmp3932;
	wire signed [31:0] w_sys_tmp3933;
	wire signed [31:0] w_sys_tmp3938;
	wire signed [31:0] w_sys_tmp3939;
	wire signed [31:0] w_sys_tmp3944;
	wire signed [31:0] w_sys_tmp3945;
	wire signed [31:0] w_sys_tmp3950;
	wire signed [31:0] w_sys_tmp3951;
	wire signed [31:0] w_sys_tmp3956;
	wire signed [31:0] w_sys_tmp3957;
	wire signed [31:0] w_sys_tmp3961;
	wire signed [31:0] w_sys_tmp3962;
	wire signed [31:0] w_sys_tmp3966;
	wire signed [31:0] w_sys_tmp3967;
	wire signed [31:0] w_sys_tmp3971;
	wire signed [31:0] w_sys_tmp3972;
	wire signed [31:0] w_sys_tmp3976;
	wire signed [31:0] w_sys_tmp3977;
	wire signed [31:0] w_sys_tmp3981;
	wire signed [31:0] w_sys_tmp3982;
	wire signed [31:0] w_sys_tmp3986;
	wire signed [31:0] w_sys_tmp3987;
	wire signed [31:0] w_sys_tmp3991;
	wire signed [31:0] w_sys_tmp3992;
	wire signed [31:0] w_sys_tmp3996;
	wire signed [31:0] w_sys_tmp3997;
	wire signed [31:0] w_sys_tmp4001;
	wire signed [31:0] w_sys_tmp4002;
	wire signed [31:0] w_sys_tmp4006;
	wire signed [31:0] w_sys_tmp4007;
	wire signed [31:0] w_sys_tmp4011;
	wire signed [31:0] w_sys_tmp4012;
	wire signed [31:0] w_sys_tmp4016;
	wire signed [31:0] w_sys_tmp4017;
	wire signed [31:0] w_sys_tmp4021;
	wire signed [31:0] w_sys_tmp4022;
	wire signed [31:0] w_sys_tmp4026;
	wire signed [31:0] w_sys_tmp4027;
	wire signed [31:0] w_sys_tmp4031;
	wire signed [31:0] w_sys_tmp4032;
	wire signed [31:0] w_sys_tmp4036;
	wire signed [31:0] w_sys_tmp4037;
	wire signed [31:0] w_sys_tmp4041;
	wire signed [31:0] w_sys_tmp4042;
	wire signed [31:0] w_sys_tmp4046;
	wire signed [31:0] w_sys_tmp4047;
	wire signed [31:0] w_sys_tmp4051;
	wire signed [31:0] w_sys_tmp4052;
	wire signed [31:0] w_sys_tmp4056;
	wire signed [31:0] w_sys_tmp4057;
	wire signed [31:0] w_sys_tmp4061;
	wire signed [31:0] w_sys_tmp4062;
	wire signed [31:0] w_sys_tmp4066;
	wire signed [31:0] w_sys_tmp4067;
	wire signed [31:0] w_sys_tmp4071;
	wire signed [31:0] w_sys_tmp4072;
	wire signed [31:0] w_sys_tmp4076;
	wire signed [31:0] w_sys_tmp4077;
	wire signed [31:0] w_sys_tmp4081;
	wire signed [31:0] w_sys_tmp4082;
	wire signed [31:0] w_sys_tmp4086;
	wire signed [31:0] w_sys_tmp4087;
	wire signed [31:0] w_sys_tmp4091;
	wire signed [31:0] w_sys_tmp4092;
	wire signed [31:0] w_sys_tmp4096;
	wire signed [31:0] w_sys_tmp4097;
	wire signed [31:0] w_sys_tmp4101;
	wire signed [31:0] w_sys_tmp4102;
	wire signed [31:0] w_sys_tmp4106;
	wire signed [31:0] w_sys_tmp4107;
	wire signed [31:0] w_sys_tmp4111;
	wire signed [31:0] w_sys_tmp4112;
	wire signed [31:0] w_sys_tmp4116;
	wire signed [31:0] w_sys_tmp4117;
	wire signed [31:0] w_sys_tmp4121;
	wire signed [31:0] w_sys_tmp4122;
	wire signed [31:0] w_sys_tmp4126;
	wire signed [31:0] w_sys_tmp4127;
	wire signed [31:0] w_sys_tmp4131;
	wire signed [31:0] w_sys_tmp4132;
	wire signed [31:0] w_sys_tmp4136;
	wire signed [31:0] w_sys_tmp4137;
	wire signed [31:0] w_sys_tmp4141;
	wire signed [31:0] w_sys_tmp4142;
	wire signed [31:0] w_sys_tmp4146;
	wire signed [31:0] w_sys_tmp4147;
	wire signed [31:0] w_sys_tmp4151;
	wire signed [31:0] w_sys_tmp4152;
	wire signed [31:0] w_sys_tmp4156;
	wire signed [31:0] w_sys_tmp4157;
	wire signed [31:0] w_sys_tmp4161;
	wire signed [31:0] w_sys_tmp4162;
	wire signed [31:0] w_sys_tmp4166;
	wire signed [31:0] w_sys_tmp4167;
	wire signed [31:0] w_sys_tmp4171;
	wire signed [31:0] w_sys_tmp4172;
	wire signed [31:0] w_sys_tmp4176;
	wire signed [31:0] w_sys_tmp4177;
	wire signed [31:0] w_sys_tmp4181;
	wire signed [31:0] w_sys_tmp4182;
	wire signed [31:0] w_sys_tmp4186;
	wire signed [31:0] w_sys_tmp4187;
	wire signed [31:0] w_sys_tmp4191;
	wire signed [31:0] w_sys_tmp4192;
	wire signed [31:0] w_sys_tmp4196;
	wire signed [31:0] w_sys_tmp4197;
	wire signed [31:0] w_sys_tmp4201;
	wire signed [31:0] w_sys_tmp4202;
	wire signed [31:0] w_sys_tmp4206;
	wire signed [31:0] w_sys_tmp4207;
	wire signed [31:0] w_sys_tmp4211;
	wire signed [31:0] w_sys_tmp4212;
	wire signed [31:0] w_sys_tmp4216;
	wire signed [31:0] w_sys_tmp4217;
	wire signed [31:0] w_sys_tmp4221;
	wire signed [31:0] w_sys_tmp4222;
	wire signed [31:0] w_sys_tmp4226;
	wire signed [31:0] w_sys_tmp4227;
	wire signed [31:0] w_sys_tmp4231;
	wire signed [31:0] w_sys_tmp4232;
	wire signed [31:0] w_sys_tmp4236;
	wire signed [31:0] w_sys_tmp4237;
	wire signed [31:0] w_sys_tmp4241;
	wire signed [31:0] w_sys_tmp4242;
	wire signed [31:0] w_sys_tmp4246;
	wire signed [31:0] w_sys_tmp4247;
	wire signed [31:0] w_sys_tmp4251;
	wire signed [31:0] w_sys_tmp4252;
	wire signed [31:0] w_sys_tmp4256;
	wire signed [31:0] w_sys_tmp4257;
	wire signed [31:0] w_sys_tmp4261;
	wire signed [31:0] w_sys_tmp4262;
	wire signed [31:0] w_sys_tmp4266;
	wire signed [31:0] w_sys_tmp4267;
	wire signed [31:0] w_sys_tmp4271;
	wire signed [31:0] w_sys_tmp4272;
	wire signed [31:0] w_sys_tmp4276;
	wire signed [31:0] w_sys_tmp4277;
	wire signed [31:0] w_sys_tmp4281;
	wire signed [31:0] w_sys_tmp4282;
	wire signed [31:0] w_sys_tmp4286;
	wire signed [31:0] w_sys_tmp4287;
	wire signed [31:0] w_sys_tmp4291;
	wire signed [31:0] w_sys_tmp4292;
	wire signed [31:0] w_sys_tmp4296;
	wire signed [31:0] w_sys_tmp4297;
	wire signed [31:0] w_sys_tmp4301;
	wire signed [31:0] w_sys_tmp4302;
	wire signed [31:0] w_sys_tmp4306;
	wire signed [31:0] w_sys_tmp4307;
	wire signed [31:0] w_sys_tmp4311;
	wire signed [31:0] w_sys_tmp4312;
	wire signed [31:0] w_sys_tmp4316;
	wire signed [31:0] w_sys_tmp4317;
	wire signed [31:0] w_sys_tmp4321;
	wire signed [31:0] w_sys_tmp4322;
	wire signed [31:0] w_sys_tmp4326;
	wire signed [31:0] w_sys_tmp4327;
	wire signed [31:0] w_sys_tmp4331;
	wire signed [31:0] w_sys_tmp4332;
	wire signed [31:0] w_sys_tmp4336;
	wire signed [31:0] w_sys_tmp4337;
	wire signed [31:0] w_sys_tmp4341;
	wire signed [31:0] w_sys_tmp4342;
	wire signed [31:0] w_sys_tmp4346;
	wire signed [31:0] w_sys_tmp4347;
	wire signed [31:0] w_sys_tmp4351;
	wire signed [31:0] w_sys_tmp4352;
	wire signed [31:0] w_sys_tmp4356;
	wire signed [31:0] w_sys_tmp4357;
	wire signed [31:0] w_sys_tmp4361;
	wire signed [31:0] w_sys_tmp4362;
	wire signed [31:0] w_sys_tmp4366;
	wire signed [31:0] w_sys_tmp4367;
	wire signed [31:0] w_sys_tmp4371;
	wire signed [31:0] w_sys_tmp4372;
	wire signed [31:0] w_sys_tmp4376;
	wire signed [31:0] w_sys_tmp4377;
	wire signed [31:0] w_sys_tmp4381;
	wire signed [31:0] w_sys_tmp4382;
	wire signed [31:0] w_sys_tmp4386;
	wire signed [31:0] w_sys_tmp4387;
	wire signed [31:0] w_sys_tmp4391;
	wire signed [31:0] w_sys_tmp4392;
	wire signed [31:0] w_sys_tmp4396;
	wire signed [31:0] w_sys_tmp4397;
	wire signed [31:0] w_sys_tmp4401;
	wire signed [31:0] w_sys_tmp4402;
	wire signed [31:0] w_sys_tmp4406;
	wire signed [31:0] w_sys_tmp4407;
	wire signed [31:0] w_sys_tmp4411;
	wire signed [31:0] w_sys_tmp4412;
	wire signed [31:0] w_sys_tmp4416;
	wire signed [31:0] w_sys_tmp4417;
	wire signed [31:0] w_sys_tmp4421;
	wire signed [31:0] w_sys_tmp4422;
	wire signed [31:0] w_sys_tmp4426;
	wire signed [31:0] w_sys_tmp4427;
	wire signed [31:0] w_sys_tmp4431;
	wire signed [31:0] w_sys_tmp4432;
	wire signed [31:0] w_sys_tmp4436;
	wire signed [31:0] w_sys_tmp4437;
	wire signed [31:0] w_sys_tmp4441;
	wire signed [31:0] w_sys_tmp4442;
	wire signed [31:0] w_sys_tmp4446;
	wire signed [31:0] w_sys_tmp4447;
	wire signed [31:0] w_sys_tmp4451;
	wire signed [31:0] w_sys_tmp4452;
	wire signed [31:0] w_sys_tmp4456;
	wire signed [31:0] w_sys_tmp4457;
	wire signed [31:0] w_sys_tmp4461;
	wire signed [31:0] w_sys_tmp4462;
	wire signed [31:0] w_sys_tmp4466;
	wire signed [31:0] w_sys_tmp4467;
	wire signed [31:0] w_sys_tmp4471;
	wire signed [31:0] w_sys_tmp4472;
	wire signed [31:0] w_sys_tmp4476;
	wire signed [31:0] w_sys_tmp4477;
	wire signed [31:0] w_sys_tmp4481;
	wire signed [31:0] w_sys_tmp4482;
	wire signed [31:0] w_sys_tmp4486;
	wire signed [31:0] w_sys_tmp4487;
	wire signed [31:0] w_sys_tmp4491;
	wire signed [31:0] w_sys_tmp4492;
	wire signed [31:0] w_sys_tmp4496;
	wire signed [31:0] w_sys_tmp4497;
	wire signed [31:0] w_sys_tmp4501;
	wire signed [31:0] w_sys_tmp4502;
	wire signed [31:0] w_sys_tmp4505;
	wire signed [31:0] w_sys_tmp4506;
	wire               w_sys_tmp4507;
	wire               w_sys_tmp4508;
	wire signed [31:0] w_sys_tmp4509;
	wire signed [31:0] w_sys_tmp4512;
	wire signed [31:0] w_sys_tmp4513;
	wire        [31:0] w_sys_tmp4514;
	wire signed [31:0] w_sys_tmp4518;
	wire signed [31:0] w_sys_tmp4519;
	wire signed [31:0] w_sys_tmp4524;
	wire signed [31:0] w_sys_tmp4525;
	wire signed [31:0] w_sys_tmp4530;
	wire signed [31:0] w_sys_tmp4531;
	wire signed [31:0] w_sys_tmp4536;
	wire signed [31:0] w_sys_tmp4537;
	wire signed [31:0] w_sys_tmp4542;
	wire signed [31:0] w_sys_tmp4543;
	wire signed [31:0] w_sys_tmp4548;
	wire signed [31:0] w_sys_tmp4549;
	wire signed [31:0] w_sys_tmp4553;
	wire signed [31:0] w_sys_tmp4554;
	wire signed [31:0] w_sys_tmp4558;
	wire signed [31:0] w_sys_tmp4559;
	wire signed [31:0] w_sys_tmp4563;
	wire signed [31:0] w_sys_tmp4564;
	wire signed [31:0] w_sys_tmp4568;
	wire signed [31:0] w_sys_tmp4569;
	wire signed [31:0] w_sys_tmp4573;
	wire signed [31:0] w_sys_tmp4574;
	wire signed [31:0] w_sys_tmp4578;
	wire signed [31:0] w_sys_tmp4579;
	wire signed [31:0] w_sys_tmp4583;
	wire signed [31:0] w_sys_tmp4584;
	wire signed [31:0] w_sys_tmp4588;
	wire signed [31:0] w_sys_tmp4589;
	wire signed [31:0] w_sys_tmp4593;
	wire signed [31:0] w_sys_tmp4594;
	wire signed [31:0] w_sys_tmp4598;
	wire signed [31:0] w_sys_tmp4599;
	wire signed [31:0] w_sys_tmp4603;
	wire signed [31:0] w_sys_tmp4604;
	wire signed [31:0] w_sys_tmp4608;
	wire signed [31:0] w_sys_tmp4609;
	wire signed [31:0] w_sys_tmp4613;
	wire signed [31:0] w_sys_tmp4614;
	wire signed [31:0] w_sys_tmp4618;
	wire signed [31:0] w_sys_tmp4619;
	wire signed [31:0] w_sys_tmp4623;
	wire signed [31:0] w_sys_tmp4624;
	wire signed [31:0] w_sys_tmp4628;
	wire signed [31:0] w_sys_tmp4629;
	wire signed [31:0] w_sys_tmp4633;
	wire signed [31:0] w_sys_tmp4634;
	wire signed [31:0] w_sys_tmp4638;
	wire signed [31:0] w_sys_tmp4639;
	wire signed [31:0] w_sys_tmp4643;
	wire signed [31:0] w_sys_tmp4644;
	wire signed [31:0] w_sys_tmp4648;
	wire signed [31:0] w_sys_tmp4649;
	wire signed [31:0] w_sys_tmp4653;
	wire signed [31:0] w_sys_tmp4654;
	wire signed [31:0] w_sys_tmp4658;
	wire signed [31:0] w_sys_tmp4659;
	wire signed [31:0] w_sys_tmp4662;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 8'h1);
	assign w_fld_T_0_addr_0 = 10'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 10'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 10'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_fld_V_3_addr_0 = 10'sh0;
	assign w_fld_V_3_datain_0 = 32'h0;
	assign w_fld_V_3_r_w_0 = 1'h0;
	assign w_fld_V_3_ce_0 = w_sys_ce;
	assign w_fld_V_3_ce_1 = w_sys_ce;
	assign w_sub19_T_addr = ( (|r_sys_processing_methodID) ? r_sub19_T_addr : 10'sh0 ) ;
	assign w_sub19_T_datain = ( (|r_sys_processing_methodID) ? r_sub19_T_datain : 32'h0 ) ;
	assign w_sub19_T_r_w = ( (|r_sys_processing_methodID) ? r_sub19_T_r_w : 1'h0 ) ;
	assign w_sub19_V_addr = ( (|r_sys_processing_methodID) ? r_sub19_V_addr : 10'sh0 ) ;
	assign w_sub19_V_datain = ( (|r_sys_processing_methodID) ? r_sub19_V_datain : 32'h0 ) ;
	assign w_sub19_V_r_w = ( (|r_sys_processing_methodID) ? r_sub19_V_r_w : 1'h0 ) ;
	assign w_sub19_U_addr = ( (|r_sys_processing_methodID) ? r_sub19_U_addr : 10'sh0 ) ;
	assign w_sub19_U_datain = ( (|r_sys_processing_methodID) ? r_sub19_U_datain : 32'h0 ) ;
	assign w_sub19_U_r_w = ( (|r_sys_processing_methodID) ? r_sub19_U_r_w : 1'h0 ) ;
	assign w_sub19_result_addr = ( (|r_sys_processing_methodID) ? r_sub19_result_addr : 10'sh0 ) ;
	assign w_sub19_result_datain = ( (|r_sys_processing_methodID) ? r_sub19_result_datain : 32'h0 ) ;
	assign w_sub19_result_r_w = ( (|r_sys_processing_methodID) ? r_sub19_result_r_w : 1'h0 ) ;
	assign w_sub09_T_addr = ( (|r_sys_processing_methodID) ? r_sub09_T_addr : 10'sh0 ) ;
	assign w_sub09_T_datain = ( (|r_sys_processing_methodID) ? r_sub09_T_datain : 32'h0 ) ;
	assign w_sub09_T_r_w = ( (|r_sys_processing_methodID) ? r_sub09_T_r_w : 1'h0 ) ;
	assign w_sub09_V_addr = ( (|r_sys_processing_methodID) ? r_sub09_V_addr : 10'sh0 ) ;
	assign w_sub09_V_datain = ( (|r_sys_processing_methodID) ? r_sub09_V_datain : 32'h0 ) ;
	assign w_sub09_V_r_w = ( (|r_sys_processing_methodID) ? r_sub09_V_r_w : 1'h0 ) ;
	assign w_sub09_U_addr = ( (|r_sys_processing_methodID) ? r_sub09_U_addr : 10'sh0 ) ;
	assign w_sub09_U_datain = ( (|r_sys_processing_methodID) ? r_sub09_U_datain : 32'h0 ) ;
	assign w_sub09_U_r_w = ( (|r_sys_processing_methodID) ? r_sub09_U_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 10'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_T_addr = ( (|r_sys_processing_methodID) ? r_sub08_T_addr : 10'sh0 ) ;
	assign w_sub08_T_datain = ( (|r_sys_processing_methodID) ? r_sub08_T_datain : 32'h0 ) ;
	assign w_sub08_T_r_w = ( (|r_sys_processing_methodID) ? r_sub08_T_r_w : 1'h0 ) ;
	assign w_sub08_V_addr = ( (|r_sys_processing_methodID) ? r_sub08_V_addr : 10'sh0 ) ;
	assign w_sub08_V_datain = ( (|r_sys_processing_methodID) ? r_sub08_V_datain : 32'h0 ) ;
	assign w_sub08_V_r_w = ( (|r_sys_processing_methodID) ? r_sub08_V_r_w : 1'h0 ) ;
	assign w_sub08_U_addr = ( (|r_sys_processing_methodID) ? r_sub08_U_addr : 10'sh0 ) ;
	assign w_sub08_U_datain = ( (|r_sys_processing_methodID) ? r_sub08_U_datain : 32'h0 ) ;
	assign w_sub08_U_r_w = ( (|r_sys_processing_methodID) ? r_sub08_U_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 10'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub24_T_addr = ( (|r_sys_processing_methodID) ? r_sub24_T_addr : 10'sh0 ) ;
	assign w_sub24_T_datain = ( (|r_sys_processing_methodID) ? r_sub24_T_datain : 32'h0 ) ;
	assign w_sub24_T_r_w = ( (|r_sys_processing_methodID) ? r_sub24_T_r_w : 1'h0 ) ;
	assign w_sub24_V_addr = ( (|r_sys_processing_methodID) ? r_sub24_V_addr : 10'sh0 ) ;
	assign w_sub24_V_datain = ( (|r_sys_processing_methodID) ? r_sub24_V_datain : 32'h0 ) ;
	assign w_sub24_V_r_w = ( (|r_sys_processing_methodID) ? r_sub24_V_r_w : 1'h0 ) ;
	assign w_sub24_U_addr = ( (|r_sys_processing_methodID) ? r_sub24_U_addr : 10'sh0 ) ;
	assign w_sub24_U_datain = ( (|r_sys_processing_methodID) ? r_sub24_U_datain : 32'h0 ) ;
	assign w_sub24_U_r_w = ( (|r_sys_processing_methodID) ? r_sub24_U_r_w : 1'h0 ) ;
	assign w_sub24_result_addr = ( (|r_sys_processing_methodID) ? r_sub24_result_addr : 10'sh0 ) ;
	assign w_sub24_result_datain = ( (|r_sys_processing_methodID) ? r_sub24_result_datain : 32'h0 ) ;
	assign w_sub24_result_r_w = ( (|r_sys_processing_methodID) ? r_sub24_result_r_w : 1'h0 ) ;
	assign w_sub22_T_addr = ( (|r_sys_processing_methodID) ? r_sub22_T_addr : 10'sh0 ) ;
	assign w_sub22_T_datain = ( (|r_sys_processing_methodID) ? r_sub22_T_datain : 32'h0 ) ;
	assign w_sub22_T_r_w = ( (|r_sys_processing_methodID) ? r_sub22_T_r_w : 1'h0 ) ;
	assign w_sub22_V_addr = ( (|r_sys_processing_methodID) ? r_sub22_V_addr : 10'sh0 ) ;
	assign w_sub22_V_datain = ( (|r_sys_processing_methodID) ? r_sub22_V_datain : 32'h0 ) ;
	assign w_sub22_V_r_w = ( (|r_sys_processing_methodID) ? r_sub22_V_r_w : 1'h0 ) ;
	assign w_sub22_U_addr = ( (|r_sys_processing_methodID) ? r_sub22_U_addr : 10'sh0 ) ;
	assign w_sub22_U_datain = ( (|r_sys_processing_methodID) ? r_sub22_U_datain : 32'h0 ) ;
	assign w_sub22_U_r_w = ( (|r_sys_processing_methodID) ? r_sub22_U_r_w : 1'h0 ) ;
	assign w_sub22_result_addr = ( (|r_sys_processing_methodID) ? r_sub22_result_addr : 10'sh0 ) ;
	assign w_sub22_result_datain = ( (|r_sys_processing_methodID) ? r_sub22_result_datain : 32'h0 ) ;
	assign w_sub22_result_r_w = ( (|r_sys_processing_methodID) ? r_sub22_result_r_w : 1'h0 ) ;
	assign w_sub23_T_addr = ( (|r_sys_processing_methodID) ? r_sub23_T_addr : 10'sh0 ) ;
	assign w_sub23_T_datain = ( (|r_sys_processing_methodID) ? r_sub23_T_datain : 32'h0 ) ;
	assign w_sub23_T_r_w = ( (|r_sys_processing_methodID) ? r_sub23_T_r_w : 1'h0 ) ;
	assign w_sub23_V_addr = ( (|r_sys_processing_methodID) ? r_sub23_V_addr : 10'sh0 ) ;
	assign w_sub23_V_datain = ( (|r_sys_processing_methodID) ? r_sub23_V_datain : 32'h0 ) ;
	assign w_sub23_V_r_w = ( (|r_sys_processing_methodID) ? r_sub23_V_r_w : 1'h0 ) ;
	assign w_sub23_U_addr = ( (|r_sys_processing_methodID) ? r_sub23_U_addr : 10'sh0 ) ;
	assign w_sub23_U_datain = ( (|r_sys_processing_methodID) ? r_sub23_U_datain : 32'h0 ) ;
	assign w_sub23_U_r_w = ( (|r_sys_processing_methodID) ? r_sub23_U_r_w : 1'h0 ) ;
	assign w_sub23_result_addr = ( (|r_sys_processing_methodID) ? r_sub23_result_addr : 10'sh0 ) ;
	assign w_sub23_result_datain = ( (|r_sys_processing_methodID) ? r_sub23_result_datain : 32'h0 ) ;
	assign w_sub23_result_r_w = ( (|r_sys_processing_methodID) ? r_sub23_result_r_w : 1'h0 ) ;
	assign w_sub12_T_addr = ( (|r_sys_processing_methodID) ? r_sub12_T_addr : 10'sh0 ) ;
	assign w_sub12_T_datain = ( (|r_sys_processing_methodID) ? r_sub12_T_datain : 32'h0 ) ;
	assign w_sub12_T_r_w = ( (|r_sys_processing_methodID) ? r_sub12_T_r_w : 1'h0 ) ;
	assign w_sub12_V_addr = ( (|r_sys_processing_methodID) ? r_sub12_V_addr : 10'sh0 ) ;
	assign w_sub12_V_datain = ( (|r_sys_processing_methodID) ? r_sub12_V_datain : 32'h0 ) ;
	assign w_sub12_V_r_w = ( (|r_sys_processing_methodID) ? r_sub12_V_r_w : 1'h0 ) ;
	assign w_sub12_U_addr = ( (|r_sys_processing_methodID) ? r_sub12_U_addr : 10'sh0 ) ;
	assign w_sub12_U_datain = ( (|r_sys_processing_methodID) ? r_sub12_U_datain : 32'h0 ) ;
	assign w_sub12_U_r_w = ( (|r_sys_processing_methodID) ? r_sub12_U_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 10'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_T_addr = ( (|r_sys_processing_methodID) ? r_sub03_T_addr : 10'sh0 ) ;
	assign w_sub03_T_datain = ( (|r_sys_processing_methodID) ? r_sub03_T_datain : 32'h0 ) ;
	assign w_sub03_T_r_w = ( (|r_sys_processing_methodID) ? r_sub03_T_r_w : 1'h0 ) ;
	assign w_sub03_V_addr = ( (|r_sys_processing_methodID) ? r_sub03_V_addr : 10'sh0 ) ;
	assign w_sub03_V_datain = ( (|r_sys_processing_methodID) ? r_sub03_V_datain : 32'h0 ) ;
	assign w_sub03_V_r_w = ( (|r_sys_processing_methodID) ? r_sub03_V_r_w : 1'h0 ) ;
	assign w_sub03_U_addr = ( (|r_sys_processing_methodID) ? r_sub03_U_addr : 10'sh0 ) ;
	assign w_sub03_U_datain = ( (|r_sys_processing_methodID) ? r_sub03_U_datain : 32'h0 ) ;
	assign w_sub03_U_r_w = ( (|r_sys_processing_methodID) ? r_sub03_U_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 10'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_T_addr = ( (|r_sys_processing_methodID) ? r_sub02_T_addr : 10'sh0 ) ;
	assign w_sub02_T_datain = ( (|r_sys_processing_methodID) ? r_sub02_T_datain : 32'h0 ) ;
	assign w_sub02_T_r_w = ( (|r_sys_processing_methodID) ? r_sub02_T_r_w : 1'h0 ) ;
	assign w_sub02_V_addr = ( (|r_sys_processing_methodID) ? r_sub02_V_addr : 10'sh0 ) ;
	assign w_sub02_V_datain = ( (|r_sys_processing_methodID) ? r_sub02_V_datain : 32'h0 ) ;
	assign w_sub02_V_r_w = ( (|r_sys_processing_methodID) ? r_sub02_V_r_w : 1'h0 ) ;
	assign w_sub02_U_addr = ( (|r_sys_processing_methodID) ? r_sub02_U_addr : 10'sh0 ) ;
	assign w_sub02_U_datain = ( (|r_sys_processing_methodID) ? r_sub02_U_datain : 32'h0 ) ;
	assign w_sub02_U_r_w = ( (|r_sys_processing_methodID) ? r_sub02_U_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 10'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_T_addr = ( (|r_sys_processing_methodID) ? r_sub11_T_addr : 10'sh0 ) ;
	assign w_sub11_T_datain = ( (|r_sys_processing_methodID) ? r_sub11_T_datain : 32'h0 ) ;
	assign w_sub11_T_r_w = ( (|r_sys_processing_methodID) ? r_sub11_T_r_w : 1'h0 ) ;
	assign w_sub11_V_addr = ( (|r_sys_processing_methodID) ? r_sub11_V_addr : 10'sh0 ) ;
	assign w_sub11_V_datain = ( (|r_sys_processing_methodID) ? r_sub11_V_datain : 32'h0 ) ;
	assign w_sub11_V_r_w = ( (|r_sys_processing_methodID) ? r_sub11_V_r_w : 1'h0 ) ;
	assign w_sub11_U_addr = ( (|r_sys_processing_methodID) ? r_sub11_U_addr : 10'sh0 ) ;
	assign w_sub11_U_datain = ( (|r_sys_processing_methodID) ? r_sub11_U_datain : 32'h0 ) ;
	assign w_sub11_U_r_w = ( (|r_sys_processing_methodID) ? r_sub11_U_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 10'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_T_addr = ( (|r_sys_processing_methodID) ? r_sub14_T_addr : 10'sh0 ) ;
	assign w_sub14_T_datain = ( (|r_sys_processing_methodID) ? r_sub14_T_datain : 32'h0 ) ;
	assign w_sub14_T_r_w = ( (|r_sys_processing_methodID) ? r_sub14_T_r_w : 1'h0 ) ;
	assign w_sub14_V_addr = ( (|r_sys_processing_methodID) ? r_sub14_V_addr : 10'sh0 ) ;
	assign w_sub14_V_datain = ( (|r_sys_processing_methodID) ? r_sub14_V_datain : 32'h0 ) ;
	assign w_sub14_V_r_w = ( (|r_sys_processing_methodID) ? r_sub14_V_r_w : 1'h0 ) ;
	assign w_sub14_U_addr = ( (|r_sys_processing_methodID) ? r_sub14_U_addr : 10'sh0 ) ;
	assign w_sub14_U_datain = ( (|r_sys_processing_methodID) ? r_sub14_U_datain : 32'h0 ) ;
	assign w_sub14_U_r_w = ( (|r_sys_processing_methodID) ? r_sub14_U_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 10'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_T_addr = ( (|r_sys_processing_methodID) ? r_sub01_T_addr : 10'sh0 ) ;
	assign w_sub01_T_datain = ( (|r_sys_processing_methodID) ? r_sub01_T_datain : 32'h0 ) ;
	assign w_sub01_T_r_w = ( (|r_sys_processing_methodID) ? r_sub01_T_r_w : 1'h0 ) ;
	assign w_sub01_V_addr = ( (|r_sys_processing_methodID) ? r_sub01_V_addr : 10'sh0 ) ;
	assign w_sub01_V_datain = ( (|r_sys_processing_methodID) ? r_sub01_V_datain : 32'h0 ) ;
	assign w_sub01_V_r_w = ( (|r_sys_processing_methodID) ? r_sub01_V_r_w : 1'h0 ) ;
	assign w_sub01_U_addr = ( (|r_sys_processing_methodID) ? r_sub01_U_addr : 10'sh0 ) ;
	assign w_sub01_U_datain = ( (|r_sys_processing_methodID) ? r_sub01_U_datain : 32'h0 ) ;
	assign w_sub01_U_r_w = ( (|r_sys_processing_methodID) ? r_sub01_U_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 10'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_T_addr = ( (|r_sys_processing_methodID) ? r_sub00_T_addr : 10'sh0 ) ;
	assign w_sub00_T_datain = ( (|r_sys_processing_methodID) ? r_sub00_T_datain : 32'h0 ) ;
	assign w_sub00_T_r_w = ( (|r_sys_processing_methodID) ? r_sub00_T_r_w : 1'h0 ) ;
	assign w_sub00_V_addr = ( (|r_sys_processing_methodID) ? r_sub00_V_addr : 10'sh0 ) ;
	assign w_sub00_V_datain = ( (|r_sys_processing_methodID) ? r_sub00_V_datain : 32'h0 ) ;
	assign w_sub00_V_r_w = ( (|r_sys_processing_methodID) ? r_sub00_V_r_w : 1'h0 ) ;
	assign w_sub00_U_addr = ( (|r_sys_processing_methodID) ? r_sub00_U_addr : 10'sh0 ) ;
	assign w_sub00_U_datain = ( (|r_sys_processing_methodID) ? r_sub00_U_datain : 32'h0 ) ;
	assign w_sub00_U_r_w = ( (|r_sys_processing_methodID) ? r_sub00_U_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 10'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub13_T_addr = ( (|r_sys_processing_methodID) ? r_sub13_T_addr : 10'sh0 ) ;
	assign w_sub13_T_datain = ( (|r_sys_processing_methodID) ? r_sub13_T_datain : 32'h0 ) ;
	assign w_sub13_T_r_w = ( (|r_sys_processing_methodID) ? r_sub13_T_r_w : 1'h0 ) ;
	assign w_sub13_V_addr = ( (|r_sys_processing_methodID) ? r_sub13_V_addr : 10'sh0 ) ;
	assign w_sub13_V_datain = ( (|r_sys_processing_methodID) ? r_sub13_V_datain : 32'h0 ) ;
	assign w_sub13_V_r_w = ( (|r_sys_processing_methodID) ? r_sub13_V_r_w : 1'h0 ) ;
	assign w_sub13_U_addr = ( (|r_sys_processing_methodID) ? r_sub13_U_addr : 10'sh0 ) ;
	assign w_sub13_U_datain = ( (|r_sys_processing_methodID) ? r_sub13_U_datain : 32'h0 ) ;
	assign w_sub13_U_r_w = ( (|r_sys_processing_methodID) ? r_sub13_U_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 10'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub07_T_addr = ( (|r_sys_processing_methodID) ? r_sub07_T_addr : 10'sh0 ) ;
	assign w_sub07_T_datain = ( (|r_sys_processing_methodID) ? r_sub07_T_datain : 32'h0 ) ;
	assign w_sub07_T_r_w = ( (|r_sys_processing_methodID) ? r_sub07_T_r_w : 1'h0 ) ;
	assign w_sub07_V_addr = ( (|r_sys_processing_methodID) ? r_sub07_V_addr : 10'sh0 ) ;
	assign w_sub07_V_datain = ( (|r_sys_processing_methodID) ? r_sub07_V_datain : 32'h0 ) ;
	assign w_sub07_V_r_w = ( (|r_sys_processing_methodID) ? r_sub07_V_r_w : 1'h0 ) ;
	assign w_sub07_U_addr = ( (|r_sys_processing_methodID) ? r_sub07_U_addr : 10'sh0 ) ;
	assign w_sub07_U_datain = ( (|r_sys_processing_methodID) ? r_sub07_U_datain : 32'h0 ) ;
	assign w_sub07_U_r_w = ( (|r_sys_processing_methodID) ? r_sub07_U_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 10'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub16_T_addr = ( (|r_sys_processing_methodID) ? r_sub16_T_addr : 10'sh0 ) ;
	assign w_sub16_T_datain = ( (|r_sys_processing_methodID) ? r_sub16_T_datain : 32'h0 ) ;
	assign w_sub16_T_r_w = ( (|r_sys_processing_methodID) ? r_sub16_T_r_w : 1'h0 ) ;
	assign w_sub16_V_addr = ( (|r_sys_processing_methodID) ? r_sub16_V_addr : 10'sh0 ) ;
	assign w_sub16_V_datain = ( (|r_sys_processing_methodID) ? r_sub16_V_datain : 32'h0 ) ;
	assign w_sub16_V_r_w = ( (|r_sys_processing_methodID) ? r_sub16_V_r_w : 1'h0 ) ;
	assign w_sub16_U_addr = ( (|r_sys_processing_methodID) ? r_sub16_U_addr : 10'sh0 ) ;
	assign w_sub16_U_datain = ( (|r_sys_processing_methodID) ? r_sub16_U_datain : 32'h0 ) ;
	assign w_sub16_U_r_w = ( (|r_sys_processing_methodID) ? r_sub16_U_r_w : 1'h0 ) ;
	assign w_sub16_result_addr = ( (|r_sys_processing_methodID) ? r_sub16_result_addr : 10'sh0 ) ;
	assign w_sub16_result_datain = ( (|r_sys_processing_methodID) ? r_sub16_result_datain : 32'h0 ) ;
	assign w_sub16_result_r_w = ( (|r_sys_processing_methodID) ? r_sub16_result_r_w : 1'h0 ) ;
	assign w_sub06_T_addr = ( (|r_sys_processing_methodID) ? r_sub06_T_addr : 10'sh0 ) ;
	assign w_sub06_T_datain = ( (|r_sys_processing_methodID) ? r_sub06_T_datain : 32'h0 ) ;
	assign w_sub06_T_r_w = ( (|r_sys_processing_methodID) ? r_sub06_T_r_w : 1'h0 ) ;
	assign w_sub06_V_addr = ( (|r_sys_processing_methodID) ? r_sub06_V_addr : 10'sh0 ) ;
	assign w_sub06_V_datain = ( (|r_sys_processing_methodID) ? r_sub06_V_datain : 32'h0 ) ;
	assign w_sub06_V_r_w = ( (|r_sys_processing_methodID) ? r_sub06_V_r_w : 1'h0 ) ;
	assign w_sub06_U_addr = ( (|r_sys_processing_methodID) ? r_sub06_U_addr : 10'sh0 ) ;
	assign w_sub06_U_datain = ( (|r_sys_processing_methodID) ? r_sub06_U_datain : 32'h0 ) ;
	assign w_sub06_U_r_w = ( (|r_sys_processing_methodID) ? r_sub06_U_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 10'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_T_addr = ( (|r_sys_processing_methodID) ? r_sub15_T_addr : 10'sh0 ) ;
	assign w_sub15_T_datain = ( (|r_sys_processing_methodID) ? r_sub15_T_datain : 32'h0 ) ;
	assign w_sub15_T_r_w = ( (|r_sys_processing_methodID) ? r_sub15_T_r_w : 1'h0 ) ;
	assign w_sub15_V_addr = ( (|r_sys_processing_methodID) ? r_sub15_V_addr : 10'sh0 ) ;
	assign w_sub15_V_datain = ( (|r_sys_processing_methodID) ? r_sub15_V_datain : 32'h0 ) ;
	assign w_sub15_V_r_w = ( (|r_sys_processing_methodID) ? r_sub15_V_r_w : 1'h0 ) ;
	assign w_sub15_U_addr = ( (|r_sys_processing_methodID) ? r_sub15_U_addr : 10'sh0 ) ;
	assign w_sub15_U_datain = ( (|r_sys_processing_methodID) ? r_sub15_U_datain : 32'h0 ) ;
	assign w_sub15_U_r_w = ( (|r_sys_processing_methodID) ? r_sub15_U_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 10'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_T_addr = ( (|r_sys_processing_methodID) ? r_sub05_T_addr : 10'sh0 ) ;
	assign w_sub05_T_datain = ( (|r_sys_processing_methodID) ? r_sub05_T_datain : 32'h0 ) ;
	assign w_sub05_T_r_w = ( (|r_sys_processing_methodID) ? r_sub05_T_r_w : 1'h0 ) ;
	assign w_sub05_V_addr = ( (|r_sys_processing_methodID) ? r_sub05_V_addr : 10'sh0 ) ;
	assign w_sub05_V_datain = ( (|r_sys_processing_methodID) ? r_sub05_V_datain : 32'h0 ) ;
	assign w_sub05_V_r_w = ( (|r_sys_processing_methodID) ? r_sub05_V_r_w : 1'h0 ) ;
	assign w_sub05_U_addr = ( (|r_sys_processing_methodID) ? r_sub05_U_addr : 10'sh0 ) ;
	assign w_sub05_U_datain = ( (|r_sys_processing_methodID) ? r_sub05_U_datain : 32'h0 ) ;
	assign w_sub05_U_r_w = ( (|r_sys_processing_methodID) ? r_sub05_U_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 10'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub18_T_addr = ( (|r_sys_processing_methodID) ? r_sub18_T_addr : 10'sh0 ) ;
	assign w_sub18_T_datain = ( (|r_sys_processing_methodID) ? r_sub18_T_datain : 32'h0 ) ;
	assign w_sub18_T_r_w = ( (|r_sys_processing_methodID) ? r_sub18_T_r_w : 1'h0 ) ;
	assign w_sub18_V_addr = ( (|r_sys_processing_methodID) ? r_sub18_V_addr : 10'sh0 ) ;
	assign w_sub18_V_datain = ( (|r_sys_processing_methodID) ? r_sub18_V_datain : 32'h0 ) ;
	assign w_sub18_V_r_w = ( (|r_sys_processing_methodID) ? r_sub18_V_r_w : 1'h0 ) ;
	assign w_sub18_U_addr = ( (|r_sys_processing_methodID) ? r_sub18_U_addr : 10'sh0 ) ;
	assign w_sub18_U_datain = ( (|r_sys_processing_methodID) ? r_sub18_U_datain : 32'h0 ) ;
	assign w_sub18_U_r_w = ( (|r_sys_processing_methodID) ? r_sub18_U_r_w : 1'h0 ) ;
	assign w_sub18_result_addr = ( (|r_sys_processing_methodID) ? r_sub18_result_addr : 10'sh0 ) ;
	assign w_sub18_result_datain = ( (|r_sys_processing_methodID) ? r_sub18_result_datain : 32'h0 ) ;
	assign w_sub18_result_r_w = ( (|r_sys_processing_methodID) ? r_sub18_result_r_w : 1'h0 ) ;
	assign w_sub04_T_addr = ( (|r_sys_processing_methodID) ? r_sub04_T_addr : 10'sh0 ) ;
	assign w_sub04_T_datain = ( (|r_sys_processing_methodID) ? r_sub04_T_datain : 32'h0 ) ;
	assign w_sub04_T_r_w = ( (|r_sys_processing_methodID) ? r_sub04_T_r_w : 1'h0 ) ;
	assign w_sub04_V_addr = ( (|r_sys_processing_methodID) ? r_sub04_V_addr : 10'sh0 ) ;
	assign w_sub04_V_datain = ( (|r_sys_processing_methodID) ? r_sub04_V_datain : 32'h0 ) ;
	assign w_sub04_V_r_w = ( (|r_sys_processing_methodID) ? r_sub04_V_r_w : 1'h0 ) ;
	assign w_sub04_U_addr = ( (|r_sys_processing_methodID) ? r_sub04_U_addr : 10'sh0 ) ;
	assign w_sub04_U_datain = ( (|r_sys_processing_methodID) ? r_sub04_U_datain : 32'h0 ) ;
	assign w_sub04_U_r_w = ( (|r_sys_processing_methodID) ? r_sub04_U_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 10'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub17_T_addr = ( (|r_sys_processing_methodID) ? r_sub17_T_addr : 10'sh0 ) ;
	assign w_sub17_T_datain = ( (|r_sys_processing_methodID) ? r_sub17_T_datain : 32'h0 ) ;
	assign w_sub17_T_r_w = ( (|r_sys_processing_methodID) ? r_sub17_T_r_w : 1'h0 ) ;
	assign w_sub17_V_addr = ( (|r_sys_processing_methodID) ? r_sub17_V_addr : 10'sh0 ) ;
	assign w_sub17_V_datain = ( (|r_sys_processing_methodID) ? r_sub17_V_datain : 32'h0 ) ;
	assign w_sub17_V_r_w = ( (|r_sys_processing_methodID) ? r_sub17_V_r_w : 1'h0 ) ;
	assign w_sub17_U_addr = ( (|r_sys_processing_methodID) ? r_sub17_U_addr : 10'sh0 ) ;
	assign w_sub17_U_datain = ( (|r_sys_processing_methodID) ? r_sub17_U_datain : 32'h0 ) ;
	assign w_sub17_U_r_w = ( (|r_sys_processing_methodID) ? r_sub17_U_r_w : 1'h0 ) ;
	assign w_sub17_result_addr = ( (|r_sys_processing_methodID) ? r_sub17_result_addr : 10'sh0 ) ;
	assign w_sub17_result_datain = ( (|r_sys_processing_methodID) ? r_sub17_result_datain : 32'h0 ) ;
	assign w_sub17_result_r_w = ( (|r_sys_processing_methodID) ? r_sub17_result_r_w : 1'h0 ) ;
	assign w_sub10_T_addr = ( (|r_sys_processing_methodID) ? r_sub10_T_addr : 10'sh0 ) ;
	assign w_sub10_T_datain = ( (|r_sys_processing_methodID) ? r_sub10_T_datain : 32'h0 ) ;
	assign w_sub10_T_r_w = ( (|r_sys_processing_methodID) ? r_sub10_T_r_w : 1'h0 ) ;
	assign w_sub10_V_addr = ( (|r_sys_processing_methodID) ? r_sub10_V_addr : 10'sh0 ) ;
	assign w_sub10_V_datain = ( (|r_sys_processing_methodID) ? r_sub10_V_datain : 32'h0 ) ;
	assign w_sub10_V_r_w = ( (|r_sys_processing_methodID) ? r_sub10_V_r_w : 1'h0 ) ;
	assign w_sub10_U_addr = ( (|r_sys_processing_methodID) ? r_sub10_U_addr : 10'sh0 ) ;
	assign w_sub10_U_datain = ( (|r_sys_processing_methodID) ? r_sub10_U_datain : 32'h0 ) ;
	assign w_sub10_U_r_w = ( (|r_sys_processing_methodID) ? r_sub10_U_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 10'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sub20_T_addr = ( (|r_sys_processing_methodID) ? r_sub20_T_addr : 10'sh0 ) ;
	assign w_sub20_T_datain = ( (|r_sys_processing_methodID) ? r_sub20_T_datain : 32'h0 ) ;
	assign w_sub20_T_r_w = ( (|r_sys_processing_methodID) ? r_sub20_T_r_w : 1'h0 ) ;
	assign w_sub20_V_addr = ( (|r_sys_processing_methodID) ? r_sub20_V_addr : 10'sh0 ) ;
	assign w_sub20_V_datain = ( (|r_sys_processing_methodID) ? r_sub20_V_datain : 32'h0 ) ;
	assign w_sub20_V_r_w = ( (|r_sys_processing_methodID) ? r_sub20_V_r_w : 1'h0 ) ;
	assign w_sub20_U_addr = ( (|r_sys_processing_methodID) ? r_sub20_U_addr : 10'sh0 ) ;
	assign w_sub20_U_datain = ( (|r_sys_processing_methodID) ? r_sub20_U_datain : 32'h0 ) ;
	assign w_sub20_U_r_w = ( (|r_sys_processing_methodID) ? r_sub20_U_r_w : 1'h0 ) ;
	assign w_sub20_result_addr = ( (|r_sys_processing_methodID) ? r_sub20_result_addr : 10'sh0 ) ;
	assign w_sub20_result_datain = ( (|r_sys_processing_methodID) ? r_sub20_result_datain : 32'h0 ) ;
	assign w_sub20_result_r_w = ( (|r_sys_processing_methodID) ? r_sub20_result_r_w : 1'h0 ) ;
	assign w_sub21_T_addr = ( (|r_sys_processing_methodID) ? r_sub21_T_addr : 10'sh0 ) ;
	assign w_sub21_T_datain = ( (|r_sys_processing_methodID) ? r_sub21_T_datain : 32'h0 ) ;
	assign w_sub21_T_r_w = ( (|r_sys_processing_methodID) ? r_sub21_T_r_w : 1'h0 ) ;
	assign w_sub21_V_addr = ( (|r_sys_processing_methodID) ? r_sub21_V_addr : 10'sh0 ) ;
	assign w_sub21_V_datain = ( (|r_sys_processing_methodID) ? r_sub21_V_datain : 32'h0 ) ;
	assign w_sub21_V_r_w = ( (|r_sys_processing_methodID) ? r_sub21_V_r_w : 1'h0 ) ;
	assign w_sub21_U_addr = ( (|r_sys_processing_methodID) ? r_sub21_U_addr : 10'sh0 ) ;
	assign w_sub21_U_datain = ( (|r_sys_processing_methodID) ? r_sub21_U_datain : 32'h0 ) ;
	assign w_sub21_U_r_w = ( (|r_sys_processing_methodID) ? r_sub21_U_r_w : 1'h0 ) ;
	assign w_sub21_result_addr = ( (|r_sys_processing_methodID) ? r_sub21_result_addr : 10'sh0 ) ;
	assign w_sub21_result_datain = ( (|r_sys_processing_methodID) ? r_sub21_result_datain : 32'h0 ) ;
	assign w_sub21_result_r_w = ( (|r_sys_processing_methodID) ? r_sub21_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh0000001e;
	assign w_sys_tmp3 = 32'sh0000001f;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'h3e088889;
	assign w_sys_tmp7 = 32'h3d088889;
	assign w_sys_tmp8 = 32'h3af5c28f;
	assign w_sys_tmp9 = 32'h3bf5c28f;
	assign w_sys_tmp10 = 32'h3ce66665;
	assign w_sys_tmp11 = 32'h3ee66665;
	assign w_sys_tmp12 = ( !w_sys_tmp13 );
	assign w_sys_tmp13 = (r_run_my_33 < r_run_k_29);
	assign w_sys_tmp14 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp15 = ( !w_sys_tmp16 );
	assign w_sys_tmp16 = (r_run_mx_32 < r_run_j_30);
	assign w_sys_tmp18 = w_ip_MultFloat_product_0;
	assign w_sys_tmp19 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp20 = (r_run_k_29 - w_sys_intOne);
	assign w_sys_tmp22 = (w_sys_tmp23 + r_run_k_29);
	assign w_sys_tmp23 = (r_run_j_30 * w_sys_tmp24);
	assign w_sys_tmp24 = 32'sh0000001f;
	assign w_sys_tmp25 = 32'h0;
	assign w_sys_tmp27 = (w_sys_tmp28 + r_run_k_29);
	assign w_sys_tmp28 = (r_run_copy2_j_47 * w_sys_tmp24);
	assign w_sys_tmp32 = (w_sys_tmp33 + r_run_k_29);
	assign w_sys_tmp33 = (r_run_copy1_j_46 * w_sys_tmp24);
	assign w_sys_tmp36 = 32'h42200000;
	assign w_sys_tmp37 = w_sys_tmp18;
	assign w_sys_tmp38 = 32'h3f800000;
	assign w_sys_tmp41 = (w_sys_tmp42 + r_run_k_29);
	assign w_sys_tmp42 = (r_run_copy0_j_45 * w_sys_tmp24);
	assign w_sys_tmp45 = (r_run_copy0_j_45 + w_sys_intOne);
	assign w_sys_tmp46 = (r_run_copy1_j_46 + w_sys_intOne);
	assign w_sys_tmp47 = (r_run_copy2_j_47 + w_sys_intOne);
	assign w_sys_tmp48 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp128 = r_sys_tmp4_float;
	assign w_sys_tmp226 = ( !w_sys_tmp227 );
	assign w_sys_tmp227 = (w_sys_tmp228 < r_run_k_29);
	assign w_sys_tmp228 = 32'sh00000008;
	assign w_sys_tmp231 = (w_sys_tmp232 + r_run_k_29);
	assign w_sys_tmp232 = 32'sh0000001f;
	assign w_sys_tmp233 = w_fld_U_2_dataout_1;
	assign w_sys_tmp239 = w_fld_V_3_dataout_1;
	assign w_sys_tmp243 = (w_sys_tmp244 + r_run_k_29);
	assign w_sys_tmp244 = 32'sh0000003e;
	assign w_sys_tmp255 = (w_sys_tmp256 + r_run_k_29);
	assign w_sys_tmp256 = 32'sh0000005d;
	assign w_sys_tmp267 = (w_sys_tmp268 + r_run_k_29);
	assign w_sys_tmp268 = 32'sh0000007c;
	assign w_sys_tmp279 = (w_sys_tmp280 + r_run_k_29);
	assign w_sys_tmp280 = 32'sh0000009b;
	assign w_sys_tmp291 = (w_sys_tmp292 + r_run_k_29);
	assign w_sys_tmp292 = 32'sh000000ba;
	assign w_sys_tmp303 = (w_sys_tmp304 + r_run_k_29);
	assign w_sys_tmp304 = 32'sh000000d9;
	assign w_sys_tmp315 = (w_sys_tmp316 + r_run_k_29);
	assign w_sys_tmp316 = 32'sh000000f8;
	assign w_sys_tmp351 = (w_sys_tmp352 + r_run_k_29);
	assign w_sys_tmp352 = 32'sh00000117;
	assign w_sys_tmp363 = (w_sys_tmp364 + r_run_k_29);
	assign w_sys_tmp364 = 32'sh00000136;
	assign w_sys_tmp375 = (w_sys_tmp376 + r_run_k_29);
	assign w_sys_tmp376 = 32'sh00000155;
	assign w_sys_tmp387 = (w_sys_tmp388 + r_run_k_29);
	assign w_sys_tmp388 = 32'sh00000174;
	assign w_sys_tmp399 = (w_sys_tmp400 + r_run_k_29);
	assign w_sys_tmp400 = 32'sh00000193;
	assign w_sys_tmp411 = (w_sys_tmp412 + r_run_k_29);
	assign w_sys_tmp412 = 32'sh000001b2;
	assign w_sys_tmp447 = (w_sys_tmp448 + r_run_k_29);
	assign w_sys_tmp448 = 32'sh000001d1;
	assign w_sys_tmp459 = (w_sys_tmp460 + r_run_k_29);
	assign w_sys_tmp460 = 32'sh000001f0;
	assign w_sys_tmp471 = (w_sys_tmp472 + r_run_k_29);
	assign w_sys_tmp472 = 32'sh0000020f;
	assign w_sys_tmp483 = (w_sys_tmp484 + r_run_k_29);
	assign w_sys_tmp484 = 32'sh0000022e;
	assign w_sys_tmp495 = (w_sys_tmp496 + r_run_k_29);
	assign w_sys_tmp496 = 32'sh0000024d;
	assign w_sys_tmp507 = (w_sys_tmp508 + r_run_k_29);
	assign w_sys_tmp508 = 32'sh0000026c;
	assign w_sys_tmp543 = (w_sys_tmp544 + r_run_k_29);
	assign w_sys_tmp544 = 32'sh0000028b;
	assign w_sys_tmp555 = (w_sys_tmp556 + r_run_k_29);
	assign w_sys_tmp556 = 32'sh000002aa;
	assign w_sys_tmp567 = (w_sys_tmp568 + r_run_k_29);
	assign w_sys_tmp568 = 32'sh000002c9;
	assign w_sys_tmp579 = (w_sys_tmp580 + r_run_k_29);
	assign w_sys_tmp580 = 32'sh000002e8;
	assign w_sys_tmp591 = (w_sys_tmp592 + r_run_k_29);
	assign w_sys_tmp592 = 32'sh00000307;
	assign w_sys_tmp603 = (w_sys_tmp604 + r_run_k_29);
	assign w_sys_tmp604 = 32'sh00000326;
	assign w_sys_tmp639 = (w_sys_tmp640 + r_run_k_29);
	assign w_sys_tmp640 = 32'sh00000345;
	assign w_sys_tmp651 = (w_sys_tmp652 + r_run_k_29);
	assign w_sys_tmp652 = 32'sh00000364;
	assign w_sys_tmp663 = (w_sys_tmp664 + r_run_k_29);
	assign w_sys_tmp664 = 32'sh00000383;
	assign w_sys_tmp675 = (w_sys_tmp676 + r_run_k_29);
	assign w_sys_tmp676 = 32'sh000003a2;
	assign w_sys_tmp687 = (w_sys_tmp688 + r_run_k_29);
	assign w_sys_tmp688 = 32'sh000003c1;
	assign w_sys_tmp699 = (w_sys_tmp700 + r_run_k_29);
	assign w_sys_tmp700 = 32'sh00000025;
	assign w_sys_tmp711 = (w_sys_tmp712 + r_run_k_29);
	assign w_sys_tmp712 = 32'sh00000044;
	assign w_sys_tmp723 = (w_sys_tmp724 + r_run_k_29);
	assign w_sys_tmp724 = 32'sh00000063;
	assign w_sys_tmp735 = (w_sys_tmp736 + r_run_k_29);
	assign w_sys_tmp736 = 32'sh00000082;
	assign w_sys_tmp747 = (w_sys_tmp748 + r_run_k_29);
	assign w_sys_tmp748 = 32'sh000000a1;
	assign w_sys_tmp759 = (w_sys_tmp760 + r_run_k_29);
	assign w_sys_tmp760 = 32'sh000000c0;
	assign w_sys_tmp771 = (w_sys_tmp772 + r_run_k_29);
	assign w_sys_tmp772 = 32'sh000000df;
	assign w_sys_tmp783 = (w_sys_tmp784 + r_run_k_29);
	assign w_sys_tmp784 = 32'sh000000fe;
	assign w_sys_tmp819 = (w_sys_tmp820 + r_run_k_29);
	assign w_sys_tmp820 = 32'sh0000011d;
	assign w_sys_tmp831 = (w_sys_tmp832 + r_run_k_29);
	assign w_sys_tmp832 = 32'sh0000013c;
	assign w_sys_tmp843 = (w_sys_tmp844 + r_run_k_29);
	assign w_sys_tmp844 = 32'sh0000015b;
	assign w_sys_tmp855 = (w_sys_tmp856 + r_run_k_29);
	assign w_sys_tmp856 = 32'sh0000017a;
	assign w_sys_tmp867 = (w_sys_tmp868 + r_run_k_29);
	assign w_sys_tmp868 = 32'sh00000199;
	assign w_sys_tmp879 = (w_sys_tmp880 + r_run_k_29);
	assign w_sys_tmp880 = 32'sh000001b8;
	assign w_sys_tmp915 = (w_sys_tmp916 + r_run_k_29);
	assign w_sys_tmp916 = 32'sh000001d7;
	assign w_sys_tmp927 = (w_sys_tmp928 + r_run_k_29);
	assign w_sys_tmp928 = 32'sh000001f6;
	assign w_sys_tmp939 = (w_sys_tmp940 + r_run_k_29);
	assign w_sys_tmp940 = 32'sh00000215;
	assign w_sys_tmp951 = (w_sys_tmp952 + r_run_k_29);
	assign w_sys_tmp952 = 32'sh00000234;
	assign w_sys_tmp963 = (w_sys_tmp964 + r_run_k_29);
	assign w_sys_tmp964 = 32'sh00000253;
	assign w_sys_tmp975 = (w_sys_tmp976 + r_run_k_29);
	assign w_sys_tmp976 = 32'sh00000272;
	assign w_sys_tmp1011 = (w_sys_tmp1012 + r_run_k_29);
	assign w_sys_tmp1012 = 32'sh00000291;
	assign w_sys_tmp1023 = (w_sys_tmp1024 + r_run_k_29);
	assign w_sys_tmp1024 = 32'sh000002b0;
	assign w_sys_tmp1035 = (w_sys_tmp1036 + r_run_k_29);
	assign w_sys_tmp1036 = 32'sh000002cf;
	assign w_sys_tmp1047 = (w_sys_tmp1048 + r_run_k_29);
	assign w_sys_tmp1048 = 32'sh000002ee;
	assign w_sys_tmp1059 = (w_sys_tmp1060 + r_run_k_29);
	assign w_sys_tmp1060 = 32'sh0000030d;
	assign w_sys_tmp1071 = (w_sys_tmp1072 + r_run_k_29);
	assign w_sys_tmp1072 = 32'sh0000032c;
	assign w_sys_tmp1107 = (w_sys_tmp1108 + r_run_k_29);
	assign w_sys_tmp1108 = 32'sh0000034b;
	assign w_sys_tmp1119 = (w_sys_tmp1120 + r_run_k_29);
	assign w_sys_tmp1120 = 32'sh0000036a;
	assign w_sys_tmp1131 = (w_sys_tmp1132 + r_run_k_29);
	assign w_sys_tmp1132 = 32'sh00000389;
	assign w_sys_tmp1143 = (w_sys_tmp1144 + r_run_k_29);
	assign w_sys_tmp1144 = 32'sh000003a8;
	assign w_sys_tmp1155 = (w_sys_tmp1156 + r_run_k_29);
	assign w_sys_tmp1156 = 32'sh000003c7;
	assign w_sys_tmp1167 = (w_sys_tmp1168 + r_run_k_29);
	assign w_sys_tmp1168 = 32'sh0000002b;
	assign w_sys_tmp1179 = (w_sys_tmp1180 + r_run_k_29);
	assign w_sys_tmp1180 = 32'sh0000004a;
	assign w_sys_tmp1191 = (w_sys_tmp1192 + r_run_k_29);
	assign w_sys_tmp1192 = 32'sh00000069;
	assign w_sys_tmp1203 = (w_sys_tmp1204 + r_run_k_29);
	assign w_sys_tmp1204 = 32'sh00000088;
	assign w_sys_tmp1215 = (w_sys_tmp1216 + r_run_k_29);
	assign w_sys_tmp1216 = 32'sh000000a7;
	assign w_sys_tmp1227 = (w_sys_tmp1228 + r_run_k_29);
	assign w_sys_tmp1228 = 32'sh000000c6;
	assign w_sys_tmp1239 = (w_sys_tmp1240 + r_run_k_29);
	assign w_sys_tmp1240 = 32'sh000000e5;
	assign w_sys_tmp1251 = (w_sys_tmp1252 + r_run_k_29);
	assign w_sys_tmp1252 = 32'sh00000104;
	assign w_sys_tmp1287 = (w_sys_tmp1288 + r_run_k_29);
	assign w_sys_tmp1288 = 32'sh00000123;
	assign w_sys_tmp1299 = (w_sys_tmp1300 + r_run_k_29);
	assign w_sys_tmp1300 = 32'sh00000142;
	assign w_sys_tmp1311 = (w_sys_tmp1312 + r_run_k_29);
	assign w_sys_tmp1312 = 32'sh00000161;
	assign w_sys_tmp1323 = (w_sys_tmp1324 + r_run_k_29);
	assign w_sys_tmp1324 = 32'sh00000180;
	assign w_sys_tmp1335 = (w_sys_tmp1336 + r_run_k_29);
	assign w_sys_tmp1336 = 32'sh0000019f;
	assign w_sys_tmp1347 = (w_sys_tmp1348 + r_run_k_29);
	assign w_sys_tmp1348 = 32'sh000001be;
	assign w_sys_tmp1383 = (w_sys_tmp1384 + r_run_k_29);
	assign w_sys_tmp1384 = 32'sh000001dd;
	assign w_sys_tmp1395 = (w_sys_tmp1396 + r_run_k_29);
	assign w_sys_tmp1396 = 32'sh000001fc;
	assign w_sys_tmp1407 = (w_sys_tmp1408 + r_run_k_29);
	assign w_sys_tmp1408 = 32'sh0000021b;
	assign w_sys_tmp1419 = (w_sys_tmp1420 + r_run_k_29);
	assign w_sys_tmp1420 = 32'sh0000023a;
	assign w_sys_tmp1431 = (w_sys_tmp1432 + r_run_k_29);
	assign w_sys_tmp1432 = 32'sh00000259;
	assign w_sys_tmp1443 = (w_sys_tmp1444 + r_run_k_29);
	assign w_sys_tmp1444 = 32'sh00000278;
	assign w_sys_tmp1479 = (w_sys_tmp1480 + r_run_k_29);
	assign w_sys_tmp1480 = 32'sh00000297;
	assign w_sys_tmp1491 = (w_sys_tmp1492 + r_run_k_29);
	assign w_sys_tmp1492 = 32'sh000002b6;
	assign w_sys_tmp1503 = (w_sys_tmp1504 + r_run_k_29);
	assign w_sys_tmp1504 = 32'sh000002d5;
	assign w_sys_tmp1515 = (w_sys_tmp1516 + r_run_k_29);
	assign w_sys_tmp1516 = 32'sh000002f4;
	assign w_sys_tmp1527 = (w_sys_tmp1528 + r_run_k_29);
	assign w_sys_tmp1528 = 32'sh00000313;
	assign w_sys_tmp1539 = (w_sys_tmp1540 + r_run_k_29);
	assign w_sys_tmp1540 = 32'sh00000332;
	assign w_sys_tmp1575 = (w_sys_tmp1576 + r_run_k_29);
	assign w_sys_tmp1576 = 32'sh00000351;
	assign w_sys_tmp1587 = (w_sys_tmp1588 + r_run_k_29);
	assign w_sys_tmp1588 = 32'sh00000370;
	assign w_sys_tmp1599 = (w_sys_tmp1600 + r_run_k_29);
	assign w_sys_tmp1600 = 32'sh0000038f;
	assign w_sys_tmp1611 = (w_sys_tmp1612 + r_run_k_29);
	assign w_sys_tmp1612 = 32'sh000003ae;
	assign w_sys_tmp1623 = (w_sys_tmp1624 + r_run_k_29);
	assign w_sys_tmp1624 = 32'sh000003cd;
	assign w_sys_tmp1635 = (w_sys_tmp1636 + r_run_k_29);
	assign w_sys_tmp1636 = 32'sh00000031;
	assign w_sys_tmp1647 = (w_sys_tmp1648 + r_run_k_29);
	assign w_sys_tmp1648 = 32'sh00000050;
	assign w_sys_tmp1659 = (w_sys_tmp1660 + r_run_k_29);
	assign w_sys_tmp1660 = 32'sh0000006f;
	assign w_sys_tmp1671 = (w_sys_tmp1672 + r_run_k_29);
	assign w_sys_tmp1672 = 32'sh0000008e;
	assign w_sys_tmp1683 = (w_sys_tmp1684 + r_run_k_29);
	assign w_sys_tmp1684 = 32'sh000000ad;
	assign w_sys_tmp1695 = (w_sys_tmp1696 + r_run_k_29);
	assign w_sys_tmp1696 = 32'sh000000cc;
	assign w_sys_tmp1707 = (w_sys_tmp1708 + r_run_k_29);
	assign w_sys_tmp1708 = 32'sh000000eb;
	assign w_sys_tmp1719 = (w_sys_tmp1720 + r_run_k_29);
	assign w_sys_tmp1720 = 32'sh0000010a;
	assign w_sys_tmp1755 = (w_sys_tmp1756 + r_run_k_29);
	assign w_sys_tmp1756 = 32'sh00000129;
	assign w_sys_tmp1767 = (w_sys_tmp1768 + r_run_k_29);
	assign w_sys_tmp1768 = 32'sh00000148;
	assign w_sys_tmp1779 = (w_sys_tmp1780 + r_run_k_29);
	assign w_sys_tmp1780 = 32'sh00000167;
	assign w_sys_tmp1791 = (w_sys_tmp1792 + r_run_k_29);
	assign w_sys_tmp1792 = 32'sh00000186;
	assign w_sys_tmp1803 = (w_sys_tmp1804 + r_run_k_29);
	assign w_sys_tmp1804 = 32'sh000001a5;
	assign w_sys_tmp1815 = (w_sys_tmp1816 + r_run_k_29);
	assign w_sys_tmp1816 = 32'sh000001c4;
	assign w_sys_tmp1851 = (w_sys_tmp1852 + r_run_k_29);
	assign w_sys_tmp1852 = 32'sh000001e3;
	assign w_sys_tmp1863 = (w_sys_tmp1864 + r_run_k_29);
	assign w_sys_tmp1864 = 32'sh00000202;
	assign w_sys_tmp1875 = (w_sys_tmp1876 + r_run_k_29);
	assign w_sys_tmp1876 = 32'sh00000221;
	assign w_sys_tmp1887 = (w_sys_tmp1888 + r_run_k_29);
	assign w_sys_tmp1888 = 32'sh00000240;
	assign w_sys_tmp1899 = (w_sys_tmp1900 + r_run_k_29);
	assign w_sys_tmp1900 = 32'sh0000025f;
	assign w_sys_tmp1911 = (w_sys_tmp1912 + r_run_k_29);
	assign w_sys_tmp1912 = 32'sh0000027e;
	assign w_sys_tmp1947 = (w_sys_tmp1948 + r_run_k_29);
	assign w_sys_tmp1948 = 32'sh0000029d;
	assign w_sys_tmp1959 = (w_sys_tmp1960 + r_run_k_29);
	assign w_sys_tmp1960 = 32'sh000002bc;
	assign w_sys_tmp1971 = (w_sys_tmp1972 + r_run_k_29);
	assign w_sys_tmp1972 = 32'sh000002db;
	assign w_sys_tmp1983 = (w_sys_tmp1984 + r_run_k_29);
	assign w_sys_tmp1984 = 32'sh000002fa;
	assign w_sys_tmp1995 = (w_sys_tmp1996 + r_run_k_29);
	assign w_sys_tmp1996 = 32'sh00000319;
	assign w_sys_tmp2007 = (w_sys_tmp2008 + r_run_k_29);
	assign w_sys_tmp2008 = 32'sh00000338;
	assign w_sys_tmp2043 = (w_sys_tmp2044 + r_run_k_29);
	assign w_sys_tmp2044 = 32'sh00000357;
	assign w_sys_tmp2055 = (w_sys_tmp2056 + r_run_k_29);
	assign w_sys_tmp2056 = 32'sh00000376;
	assign w_sys_tmp2067 = (w_sys_tmp2068 + r_run_k_29);
	assign w_sys_tmp2068 = 32'sh00000395;
	assign w_sys_tmp2079 = (w_sys_tmp2080 + r_run_k_29);
	assign w_sys_tmp2080 = 32'sh000003b4;
	assign w_sys_tmp2091 = (w_sys_tmp2092 + r_run_k_29);
	assign w_sys_tmp2092 = 32'sh000003d3;
	assign w_sys_tmp2102 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp2103 = 32'sh00000019;
	assign w_sys_tmp2104 = ( !w_sys_tmp2105 );
	assign w_sys_tmp2105 = (w_sys_tmp2106 < r_run_k_29);
	assign w_sys_tmp2106 = 32'sh0000001f;
	assign w_sys_tmp2109 = (w_sys_tmp2110 + r_run_k_29);
	assign w_sys_tmp2110 = 32'sh0000001f;
	assign w_sys_tmp2111 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2117 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2121 = (w_sys_tmp2122 + r_run_k_29);
	assign w_sys_tmp2122 = 32'sh0000003e;
	assign w_sys_tmp2133 = (w_sys_tmp2134 + r_run_k_29);
	assign w_sys_tmp2134 = 32'sh0000005d;
	assign w_sys_tmp2145 = (w_sys_tmp2146 + r_run_k_29);
	assign w_sys_tmp2146 = 32'sh0000007c;
	assign w_sys_tmp2157 = (w_sys_tmp2158 + r_run_k_29);
	assign w_sys_tmp2158 = 32'sh0000009b;
	assign w_sys_tmp2169 = (w_sys_tmp2170 + r_run_k_29);
	assign w_sys_tmp2170 = 32'sh000000ba;
	assign w_sys_tmp2181 = (w_sys_tmp2182 + r_run_k_29);
	assign w_sys_tmp2182 = 32'sh000000d9;
	assign w_sys_tmp2193 = (w_sys_tmp2194 + r_run_k_29);
	assign w_sys_tmp2194 = 32'sh000000f8;
	assign w_sys_tmp2229 = (w_sys_tmp2230 + r_run_k_29);
	assign w_sys_tmp2230 = 32'sh00000117;
	assign w_sys_tmp2241 = (w_sys_tmp2242 + r_run_k_29);
	assign w_sys_tmp2242 = 32'sh00000136;
	assign w_sys_tmp2253 = (w_sys_tmp2254 + r_run_k_29);
	assign w_sys_tmp2254 = 32'sh00000155;
	assign w_sys_tmp2265 = (w_sys_tmp2266 + r_run_k_29);
	assign w_sys_tmp2266 = 32'sh00000174;
	assign w_sys_tmp2277 = (w_sys_tmp2278 + r_run_k_29);
	assign w_sys_tmp2278 = 32'sh00000193;
	assign w_sys_tmp2289 = (w_sys_tmp2290 + r_run_k_29);
	assign w_sys_tmp2290 = 32'sh000001b2;
	assign w_sys_tmp2325 = (w_sys_tmp2326 + r_run_k_29);
	assign w_sys_tmp2326 = 32'sh000001d1;
	assign w_sys_tmp2337 = (w_sys_tmp2338 + r_run_k_29);
	assign w_sys_tmp2338 = 32'sh000001f0;
	assign w_sys_tmp2349 = (w_sys_tmp2350 + r_run_k_29);
	assign w_sys_tmp2350 = 32'sh0000020f;
	assign w_sys_tmp2361 = (w_sys_tmp2362 + r_run_k_29);
	assign w_sys_tmp2362 = 32'sh0000022e;
	assign w_sys_tmp2373 = (w_sys_tmp2374 + r_run_k_29);
	assign w_sys_tmp2374 = 32'sh0000024d;
	assign w_sys_tmp2385 = (w_sys_tmp2386 + r_run_k_29);
	assign w_sys_tmp2386 = 32'sh0000026c;
	assign w_sys_tmp2421 = (w_sys_tmp2422 + r_run_k_29);
	assign w_sys_tmp2422 = 32'sh0000028b;
	assign w_sys_tmp2433 = (w_sys_tmp2434 + r_run_k_29);
	assign w_sys_tmp2434 = 32'sh000002aa;
	assign w_sys_tmp2445 = (w_sys_tmp2446 + r_run_k_29);
	assign w_sys_tmp2446 = 32'sh000002c9;
	assign w_sys_tmp2457 = (w_sys_tmp2458 + r_run_k_29);
	assign w_sys_tmp2458 = 32'sh000002e8;
	assign w_sys_tmp2469 = (w_sys_tmp2470 + r_run_k_29);
	assign w_sys_tmp2470 = 32'sh00000307;
	assign w_sys_tmp2481 = (w_sys_tmp2482 + r_run_k_29);
	assign w_sys_tmp2482 = 32'sh00000326;
	assign w_sys_tmp2517 = (w_sys_tmp2518 + r_run_k_29);
	assign w_sys_tmp2518 = 32'sh00000345;
	assign w_sys_tmp2529 = (w_sys_tmp2530 + r_run_k_29);
	assign w_sys_tmp2530 = 32'sh00000364;
	assign w_sys_tmp2541 = (w_sys_tmp2542 + r_run_k_29);
	assign w_sys_tmp2542 = 32'sh00000383;
	assign w_sys_tmp2553 = (w_sys_tmp2554 + r_run_k_29);
	assign w_sys_tmp2554 = 32'sh000003a2;
	assign w_sys_tmp2565 = (w_sys_tmp2566 + r_run_k_29);
	assign w_sys_tmp2566 = 32'sh000003c1;
	assign w_sys_tmp2576 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp2577 = ( !w_sys_tmp2578 );
	assign w_sys_tmp2578 = (r_run_nlast_44 < r_run_n_31);
	assign w_sys_tmp2579 = (r_run_n_31 + w_sys_intOne);
	assign w_sys_tmp2580 = ( !w_sys_tmp2581 );
	assign w_sys_tmp2581 = (r_run_my_33 < r_run_k_29);
	assign w_sys_tmp2584 = (w_sys_tmp2585 + r_run_k_29);
	assign w_sys_tmp2585 = 32'sh0000001f;
	assign w_sys_tmp2586 = 32'h0;
	assign w_sys_tmp2588 = (w_sys_tmp2589 + r_run_k_29);
	assign w_sys_tmp2589 = (r_run_mx_32 * w_sys_tmp2585);
	assign w_sys_tmp2591 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2592 = (w_sys_tmp2593 + r_run_k_29);
	assign w_sys_tmp2593 = (w_sys_tmp2594 * w_sys_tmp2585);
	assign w_sys_tmp2594 = (r_run_mx_32 - w_sys_intOne);
	assign w_sys_tmp2596 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp2597 = ( !w_sys_tmp2598 );
	assign w_sys_tmp2598 = (r_run_mx_32 < r_run_j_30);
	assign w_sys_tmp2601 = (w_sys_tmp2602 + w_sys_intOne);
	assign w_sys_tmp2602 = (r_run_j_30 * w_sys_tmp2603);
	assign w_sys_tmp2603 = 32'sh0000001f;
	assign w_sys_tmp2604 = 32'h0;
	assign w_sys_tmp2606 = (w_sys_tmp2607 + r_run_my_33);
	assign w_sys_tmp2607 = (r_run_copy0_j_48 * w_sys_tmp2603);
	assign w_sys_tmp2610 = (r_run_copy0_j_48 + w_sys_intOne);
	assign w_sys_tmp2611 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp2684 = w_ip_DivInt_quotient_0;
	assign w_sys_tmp2685 = 32'sh00000004;
	assign w_sys_tmp2686 = ( !w_sys_tmp2687 );
	assign w_sys_tmp2687 = (w_sys_tmp2688 < r_run_j_30);
	assign w_sys_tmp2688 = w_ip_DivInt_quotient_1;
	assign w_sys_tmp2689 = 32'sh00000002;
	assign w_sys_tmp2692 = (w_sys_tmp2693 + w_sys_intOne);
	assign w_sys_tmp2693 = (r_run_j_30 * w_sys_tmp2694);
	assign w_sys_tmp2694 = 32'sh0000001f;
	assign w_sys_tmp2695 = 32'h3f800000;
	assign w_sys_tmp2696 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp2733 = ( !w_sys_tmp2734 );
	assign w_sys_tmp2734 = (w_sys_tmp2735 < r_run_k_29);
	assign w_sys_tmp2735 = 32'sh00000008;
	assign w_sys_tmp2738 = (w_sys_tmp2739 + r_run_k_29);
	assign w_sys_tmp2739 = 32'sh0000001f;
	assign w_sys_tmp2740 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2744 = (w_sys_tmp2745 + r_run_k_29);
	assign w_sys_tmp2745 = 32'sh0000003e;
	assign w_sys_tmp2750 = (w_sys_tmp2751 + r_run_k_29);
	assign w_sys_tmp2751 = 32'sh0000005d;
	assign w_sys_tmp2756 = (w_sys_tmp2757 + r_run_k_29);
	assign w_sys_tmp2757 = 32'sh0000007c;
	assign w_sys_tmp2762 = (w_sys_tmp2763 + r_run_k_29);
	assign w_sys_tmp2763 = 32'sh0000009b;
	assign w_sys_tmp2768 = (w_sys_tmp2769 + r_run_k_29);
	assign w_sys_tmp2769 = 32'sh000000ba;
	assign w_sys_tmp2774 = (w_sys_tmp2775 + r_run_k_29);
	assign w_sys_tmp2775 = 32'sh000000d9;
	assign w_sys_tmp2780 = (w_sys_tmp2781 + r_run_k_29);
	assign w_sys_tmp2781 = 32'sh000000f8;
	assign w_sys_tmp2798 = (w_sys_tmp2799 + r_run_k_29);
	assign w_sys_tmp2799 = 32'sh00000117;
	assign w_sys_tmp2804 = (w_sys_tmp2805 + r_run_k_29);
	assign w_sys_tmp2805 = 32'sh00000136;
	assign w_sys_tmp2810 = (w_sys_tmp2811 + r_run_k_29);
	assign w_sys_tmp2811 = 32'sh00000155;
	assign w_sys_tmp2816 = (w_sys_tmp2817 + r_run_k_29);
	assign w_sys_tmp2817 = 32'sh00000174;
	assign w_sys_tmp2822 = (w_sys_tmp2823 + r_run_k_29);
	assign w_sys_tmp2823 = 32'sh00000193;
	assign w_sys_tmp2828 = (w_sys_tmp2829 + r_run_k_29);
	assign w_sys_tmp2829 = 32'sh000001b2;
	assign w_sys_tmp2846 = (w_sys_tmp2847 + r_run_k_29);
	assign w_sys_tmp2847 = 32'sh000001d1;
	assign w_sys_tmp2852 = (w_sys_tmp2853 + r_run_k_29);
	assign w_sys_tmp2853 = 32'sh000001f0;
	assign w_sys_tmp2858 = (w_sys_tmp2859 + r_run_k_29);
	assign w_sys_tmp2859 = 32'sh0000020f;
	assign w_sys_tmp2864 = (w_sys_tmp2865 + r_run_k_29);
	assign w_sys_tmp2865 = 32'sh0000022e;
	assign w_sys_tmp2870 = (w_sys_tmp2871 + r_run_k_29);
	assign w_sys_tmp2871 = 32'sh0000024d;
	assign w_sys_tmp2876 = (w_sys_tmp2877 + r_run_k_29);
	assign w_sys_tmp2877 = 32'sh0000026c;
	assign w_sys_tmp2894 = (w_sys_tmp2895 + r_run_k_29);
	assign w_sys_tmp2895 = 32'sh0000028b;
	assign w_sys_tmp2900 = (w_sys_tmp2901 + r_run_k_29);
	assign w_sys_tmp2901 = 32'sh000002aa;
	assign w_sys_tmp2906 = (w_sys_tmp2907 + r_run_k_29);
	assign w_sys_tmp2907 = 32'sh000002c9;
	assign w_sys_tmp2912 = (w_sys_tmp2913 + r_run_k_29);
	assign w_sys_tmp2913 = 32'sh000002e8;
	assign w_sys_tmp2918 = (w_sys_tmp2919 + r_run_k_29);
	assign w_sys_tmp2919 = 32'sh00000307;
	assign w_sys_tmp2924 = (w_sys_tmp2925 + r_run_k_29);
	assign w_sys_tmp2925 = 32'sh00000326;
	assign w_sys_tmp2942 = (w_sys_tmp2943 + r_run_k_29);
	assign w_sys_tmp2943 = 32'sh00000345;
	assign w_sys_tmp2948 = (w_sys_tmp2949 + r_run_k_29);
	assign w_sys_tmp2949 = 32'sh00000364;
	assign w_sys_tmp2954 = (w_sys_tmp2955 + r_run_k_29);
	assign w_sys_tmp2955 = 32'sh00000383;
	assign w_sys_tmp2960 = (w_sys_tmp2961 + r_run_k_29);
	assign w_sys_tmp2961 = 32'sh000003a2;
	assign w_sys_tmp2966 = (w_sys_tmp2967 + r_run_k_29);
	assign w_sys_tmp2967 = 32'sh000003c1;
	assign w_sys_tmp2972 = (w_sys_tmp2973 + r_run_k_29);
	assign w_sys_tmp2973 = 32'sh00000025;
	assign w_sys_tmp2978 = (w_sys_tmp2979 + r_run_k_29);
	assign w_sys_tmp2979 = 32'sh00000044;
	assign w_sys_tmp2984 = (w_sys_tmp2985 + r_run_k_29);
	assign w_sys_tmp2985 = 32'sh00000063;
	assign w_sys_tmp2990 = (w_sys_tmp2991 + r_run_k_29);
	assign w_sys_tmp2991 = 32'sh00000082;
	assign w_sys_tmp2996 = (w_sys_tmp2997 + r_run_k_29);
	assign w_sys_tmp2997 = 32'sh000000a1;
	assign w_sys_tmp3002 = (w_sys_tmp3003 + r_run_k_29);
	assign w_sys_tmp3003 = 32'sh000000c0;
	assign w_sys_tmp3008 = (w_sys_tmp3009 + r_run_k_29);
	assign w_sys_tmp3009 = 32'sh000000df;
	assign w_sys_tmp3014 = (w_sys_tmp3015 + r_run_k_29);
	assign w_sys_tmp3015 = 32'sh000000fe;
	assign w_sys_tmp3032 = (w_sys_tmp3033 + r_run_k_29);
	assign w_sys_tmp3033 = 32'sh0000011d;
	assign w_sys_tmp3038 = (w_sys_tmp3039 + r_run_k_29);
	assign w_sys_tmp3039 = 32'sh0000013c;
	assign w_sys_tmp3044 = (w_sys_tmp3045 + r_run_k_29);
	assign w_sys_tmp3045 = 32'sh0000015b;
	assign w_sys_tmp3050 = (w_sys_tmp3051 + r_run_k_29);
	assign w_sys_tmp3051 = 32'sh0000017a;
	assign w_sys_tmp3056 = (w_sys_tmp3057 + r_run_k_29);
	assign w_sys_tmp3057 = 32'sh00000199;
	assign w_sys_tmp3062 = (w_sys_tmp3063 + r_run_k_29);
	assign w_sys_tmp3063 = 32'sh000001b8;
	assign w_sys_tmp3080 = (w_sys_tmp3081 + r_run_k_29);
	assign w_sys_tmp3081 = 32'sh000001d7;
	assign w_sys_tmp3086 = (w_sys_tmp3087 + r_run_k_29);
	assign w_sys_tmp3087 = 32'sh000001f6;
	assign w_sys_tmp3092 = (w_sys_tmp3093 + r_run_k_29);
	assign w_sys_tmp3093 = 32'sh00000215;
	assign w_sys_tmp3098 = (w_sys_tmp3099 + r_run_k_29);
	assign w_sys_tmp3099 = 32'sh00000234;
	assign w_sys_tmp3104 = (w_sys_tmp3105 + r_run_k_29);
	assign w_sys_tmp3105 = 32'sh00000253;
	assign w_sys_tmp3110 = (w_sys_tmp3111 + r_run_k_29);
	assign w_sys_tmp3111 = 32'sh00000272;
	assign w_sys_tmp3128 = (w_sys_tmp3129 + r_run_k_29);
	assign w_sys_tmp3129 = 32'sh00000291;
	assign w_sys_tmp3134 = (w_sys_tmp3135 + r_run_k_29);
	assign w_sys_tmp3135 = 32'sh000002b0;
	assign w_sys_tmp3140 = (w_sys_tmp3141 + r_run_k_29);
	assign w_sys_tmp3141 = 32'sh000002cf;
	assign w_sys_tmp3146 = (w_sys_tmp3147 + r_run_k_29);
	assign w_sys_tmp3147 = 32'sh000002ee;
	assign w_sys_tmp3152 = (w_sys_tmp3153 + r_run_k_29);
	assign w_sys_tmp3153 = 32'sh0000030d;
	assign w_sys_tmp3158 = (w_sys_tmp3159 + r_run_k_29);
	assign w_sys_tmp3159 = 32'sh0000032c;
	assign w_sys_tmp3176 = (w_sys_tmp3177 + r_run_k_29);
	assign w_sys_tmp3177 = 32'sh0000034b;
	assign w_sys_tmp3182 = (w_sys_tmp3183 + r_run_k_29);
	assign w_sys_tmp3183 = 32'sh0000036a;
	assign w_sys_tmp3188 = (w_sys_tmp3189 + r_run_k_29);
	assign w_sys_tmp3189 = 32'sh00000389;
	assign w_sys_tmp3194 = (w_sys_tmp3195 + r_run_k_29);
	assign w_sys_tmp3195 = 32'sh000003a8;
	assign w_sys_tmp3200 = (w_sys_tmp3201 + r_run_k_29);
	assign w_sys_tmp3201 = 32'sh000003c7;
	assign w_sys_tmp3206 = (w_sys_tmp3207 + r_run_k_29);
	assign w_sys_tmp3207 = 32'sh0000002b;
	assign w_sys_tmp3212 = (w_sys_tmp3213 + r_run_k_29);
	assign w_sys_tmp3213 = 32'sh0000004a;
	assign w_sys_tmp3218 = (w_sys_tmp3219 + r_run_k_29);
	assign w_sys_tmp3219 = 32'sh00000069;
	assign w_sys_tmp3224 = (w_sys_tmp3225 + r_run_k_29);
	assign w_sys_tmp3225 = 32'sh00000088;
	assign w_sys_tmp3230 = (w_sys_tmp3231 + r_run_k_29);
	assign w_sys_tmp3231 = 32'sh000000a7;
	assign w_sys_tmp3236 = (w_sys_tmp3237 + r_run_k_29);
	assign w_sys_tmp3237 = 32'sh000000c6;
	assign w_sys_tmp3242 = (w_sys_tmp3243 + r_run_k_29);
	assign w_sys_tmp3243 = 32'sh000000e5;
	assign w_sys_tmp3248 = (w_sys_tmp3249 + r_run_k_29);
	assign w_sys_tmp3249 = 32'sh00000104;
	assign w_sys_tmp3266 = (w_sys_tmp3267 + r_run_k_29);
	assign w_sys_tmp3267 = 32'sh00000123;
	assign w_sys_tmp3272 = (w_sys_tmp3273 + r_run_k_29);
	assign w_sys_tmp3273 = 32'sh00000142;
	assign w_sys_tmp3278 = (w_sys_tmp3279 + r_run_k_29);
	assign w_sys_tmp3279 = 32'sh00000161;
	assign w_sys_tmp3284 = (w_sys_tmp3285 + r_run_k_29);
	assign w_sys_tmp3285 = 32'sh00000180;
	assign w_sys_tmp3290 = (w_sys_tmp3291 + r_run_k_29);
	assign w_sys_tmp3291 = 32'sh0000019f;
	assign w_sys_tmp3296 = (w_sys_tmp3297 + r_run_k_29);
	assign w_sys_tmp3297 = 32'sh000001be;
	assign w_sys_tmp3314 = (w_sys_tmp3315 + r_run_k_29);
	assign w_sys_tmp3315 = 32'sh000001dd;
	assign w_sys_tmp3320 = (w_sys_tmp3321 + r_run_k_29);
	assign w_sys_tmp3321 = 32'sh000001fc;
	assign w_sys_tmp3326 = (w_sys_tmp3327 + r_run_k_29);
	assign w_sys_tmp3327 = 32'sh0000021b;
	assign w_sys_tmp3332 = (w_sys_tmp3333 + r_run_k_29);
	assign w_sys_tmp3333 = 32'sh0000023a;
	assign w_sys_tmp3338 = (w_sys_tmp3339 + r_run_k_29);
	assign w_sys_tmp3339 = 32'sh00000259;
	assign w_sys_tmp3344 = (w_sys_tmp3345 + r_run_k_29);
	assign w_sys_tmp3345 = 32'sh00000278;
	assign w_sys_tmp3362 = (w_sys_tmp3363 + r_run_k_29);
	assign w_sys_tmp3363 = 32'sh00000297;
	assign w_sys_tmp3368 = (w_sys_tmp3369 + r_run_k_29);
	assign w_sys_tmp3369 = 32'sh000002b6;
	assign w_sys_tmp3374 = (w_sys_tmp3375 + r_run_k_29);
	assign w_sys_tmp3375 = 32'sh000002d5;
	assign w_sys_tmp3380 = (w_sys_tmp3381 + r_run_k_29);
	assign w_sys_tmp3381 = 32'sh000002f4;
	assign w_sys_tmp3386 = (w_sys_tmp3387 + r_run_k_29);
	assign w_sys_tmp3387 = 32'sh00000313;
	assign w_sys_tmp3392 = (w_sys_tmp3393 + r_run_k_29);
	assign w_sys_tmp3393 = 32'sh00000332;
	assign w_sys_tmp3410 = (w_sys_tmp3411 + r_run_k_29);
	assign w_sys_tmp3411 = 32'sh00000351;
	assign w_sys_tmp3416 = (w_sys_tmp3417 + r_run_k_29);
	assign w_sys_tmp3417 = 32'sh00000370;
	assign w_sys_tmp3422 = (w_sys_tmp3423 + r_run_k_29);
	assign w_sys_tmp3423 = 32'sh0000038f;
	assign w_sys_tmp3428 = (w_sys_tmp3429 + r_run_k_29);
	assign w_sys_tmp3429 = 32'sh000003ae;
	assign w_sys_tmp3434 = (w_sys_tmp3435 + r_run_k_29);
	assign w_sys_tmp3435 = 32'sh000003cd;
	assign w_sys_tmp3440 = (w_sys_tmp3441 + r_run_k_29);
	assign w_sys_tmp3441 = 32'sh00000031;
	assign w_sys_tmp3446 = (w_sys_tmp3447 + r_run_k_29);
	assign w_sys_tmp3447 = 32'sh00000050;
	assign w_sys_tmp3452 = (w_sys_tmp3453 + r_run_k_29);
	assign w_sys_tmp3453 = 32'sh0000006f;
	assign w_sys_tmp3458 = (w_sys_tmp3459 + r_run_k_29);
	assign w_sys_tmp3459 = 32'sh0000008e;
	assign w_sys_tmp3464 = (w_sys_tmp3465 + r_run_k_29);
	assign w_sys_tmp3465 = 32'sh000000ad;
	assign w_sys_tmp3470 = (w_sys_tmp3471 + r_run_k_29);
	assign w_sys_tmp3471 = 32'sh000000cc;
	assign w_sys_tmp3476 = (w_sys_tmp3477 + r_run_k_29);
	assign w_sys_tmp3477 = 32'sh000000eb;
	assign w_sys_tmp3482 = (w_sys_tmp3483 + r_run_k_29);
	assign w_sys_tmp3483 = 32'sh0000010a;
	assign w_sys_tmp3500 = (w_sys_tmp3501 + r_run_k_29);
	assign w_sys_tmp3501 = 32'sh00000129;
	assign w_sys_tmp3506 = (w_sys_tmp3507 + r_run_k_29);
	assign w_sys_tmp3507 = 32'sh00000148;
	assign w_sys_tmp3512 = (w_sys_tmp3513 + r_run_k_29);
	assign w_sys_tmp3513 = 32'sh00000167;
	assign w_sys_tmp3518 = (w_sys_tmp3519 + r_run_k_29);
	assign w_sys_tmp3519 = 32'sh00000186;
	assign w_sys_tmp3524 = (w_sys_tmp3525 + r_run_k_29);
	assign w_sys_tmp3525 = 32'sh000001a5;
	assign w_sys_tmp3530 = (w_sys_tmp3531 + r_run_k_29);
	assign w_sys_tmp3531 = 32'sh000001c4;
	assign w_sys_tmp3548 = (w_sys_tmp3549 + r_run_k_29);
	assign w_sys_tmp3549 = 32'sh000001e3;
	assign w_sys_tmp3554 = (w_sys_tmp3555 + r_run_k_29);
	assign w_sys_tmp3555 = 32'sh00000202;
	assign w_sys_tmp3560 = (w_sys_tmp3561 + r_run_k_29);
	assign w_sys_tmp3561 = 32'sh00000221;
	assign w_sys_tmp3566 = (w_sys_tmp3567 + r_run_k_29);
	assign w_sys_tmp3567 = 32'sh00000240;
	assign w_sys_tmp3572 = (w_sys_tmp3573 + r_run_k_29);
	assign w_sys_tmp3573 = 32'sh0000025f;
	assign w_sys_tmp3578 = (w_sys_tmp3579 + r_run_k_29);
	assign w_sys_tmp3579 = 32'sh0000027e;
	assign w_sys_tmp3596 = (w_sys_tmp3597 + r_run_k_29);
	assign w_sys_tmp3597 = 32'sh0000029d;
	assign w_sys_tmp3602 = (w_sys_tmp3603 + r_run_k_29);
	assign w_sys_tmp3603 = 32'sh000002bc;
	assign w_sys_tmp3608 = (w_sys_tmp3609 + r_run_k_29);
	assign w_sys_tmp3609 = 32'sh000002db;
	assign w_sys_tmp3614 = (w_sys_tmp3615 + r_run_k_29);
	assign w_sys_tmp3615 = 32'sh000002fa;
	assign w_sys_tmp3620 = (w_sys_tmp3621 + r_run_k_29);
	assign w_sys_tmp3621 = 32'sh00000319;
	assign w_sys_tmp3626 = (w_sys_tmp3627 + r_run_k_29);
	assign w_sys_tmp3627 = 32'sh00000338;
	assign w_sys_tmp3644 = (w_sys_tmp3645 + r_run_k_29);
	assign w_sys_tmp3645 = 32'sh00000357;
	assign w_sys_tmp3650 = (w_sys_tmp3651 + r_run_k_29);
	assign w_sys_tmp3651 = 32'sh00000376;
	assign w_sys_tmp3656 = (w_sys_tmp3657 + r_run_k_29);
	assign w_sys_tmp3657 = 32'sh00000395;
	assign w_sys_tmp3662 = (w_sys_tmp3663 + r_run_k_29);
	assign w_sys_tmp3663 = 32'sh000003b4;
	assign w_sys_tmp3668 = (w_sys_tmp3669 + r_run_k_29);
	assign w_sys_tmp3669 = 32'sh000003d3;
	assign w_sys_tmp3673 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp3674 = 32'sh00000019;
	assign w_sys_tmp3675 = ( !w_sys_tmp3676 );
	assign w_sys_tmp3676 = (w_sys_tmp3677 < r_run_k_29);
	assign w_sys_tmp3677 = 32'sh0000001f;
	assign w_sys_tmp3680 = (w_sys_tmp3681 + r_run_k_29);
	assign w_sys_tmp3681 = 32'sh0000001f;
	assign w_sys_tmp3682 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3686 = (w_sys_tmp3687 + r_run_k_29);
	assign w_sys_tmp3687 = 32'sh0000003e;
	assign w_sys_tmp3692 = (w_sys_tmp3693 + r_run_k_29);
	assign w_sys_tmp3693 = 32'sh0000005d;
	assign w_sys_tmp3698 = (w_sys_tmp3699 + r_run_k_29);
	assign w_sys_tmp3699 = 32'sh0000007c;
	assign w_sys_tmp3704 = (w_sys_tmp3705 + r_run_k_29);
	assign w_sys_tmp3705 = 32'sh0000009b;
	assign w_sys_tmp3710 = (w_sys_tmp3711 + r_run_k_29);
	assign w_sys_tmp3711 = 32'sh000000ba;
	assign w_sys_tmp3716 = (w_sys_tmp3717 + r_run_k_29);
	assign w_sys_tmp3717 = 32'sh000000d9;
	assign w_sys_tmp3722 = (w_sys_tmp3723 + r_run_k_29);
	assign w_sys_tmp3723 = 32'sh000000f8;
	assign w_sys_tmp3740 = (w_sys_tmp3741 + r_run_k_29);
	assign w_sys_tmp3741 = 32'sh00000117;
	assign w_sys_tmp3746 = (w_sys_tmp3747 + r_run_k_29);
	assign w_sys_tmp3747 = 32'sh00000136;
	assign w_sys_tmp3752 = (w_sys_tmp3753 + r_run_k_29);
	assign w_sys_tmp3753 = 32'sh00000155;
	assign w_sys_tmp3758 = (w_sys_tmp3759 + r_run_k_29);
	assign w_sys_tmp3759 = 32'sh00000174;
	assign w_sys_tmp3764 = (w_sys_tmp3765 + r_run_k_29);
	assign w_sys_tmp3765 = 32'sh00000193;
	assign w_sys_tmp3770 = (w_sys_tmp3771 + r_run_k_29);
	assign w_sys_tmp3771 = 32'sh000001b2;
	assign w_sys_tmp3788 = (w_sys_tmp3789 + r_run_k_29);
	assign w_sys_tmp3789 = 32'sh000001d1;
	assign w_sys_tmp3794 = (w_sys_tmp3795 + r_run_k_29);
	assign w_sys_tmp3795 = 32'sh000001f0;
	assign w_sys_tmp3800 = (w_sys_tmp3801 + r_run_k_29);
	assign w_sys_tmp3801 = 32'sh0000020f;
	assign w_sys_tmp3806 = (w_sys_tmp3807 + r_run_k_29);
	assign w_sys_tmp3807 = 32'sh0000022e;
	assign w_sys_tmp3812 = (w_sys_tmp3813 + r_run_k_29);
	assign w_sys_tmp3813 = 32'sh0000024d;
	assign w_sys_tmp3818 = (w_sys_tmp3819 + r_run_k_29);
	assign w_sys_tmp3819 = 32'sh0000026c;
	assign w_sys_tmp3836 = (w_sys_tmp3837 + r_run_k_29);
	assign w_sys_tmp3837 = 32'sh0000028b;
	assign w_sys_tmp3842 = (w_sys_tmp3843 + r_run_k_29);
	assign w_sys_tmp3843 = 32'sh000002aa;
	assign w_sys_tmp3848 = (w_sys_tmp3849 + r_run_k_29);
	assign w_sys_tmp3849 = 32'sh000002c9;
	assign w_sys_tmp3854 = (w_sys_tmp3855 + r_run_k_29);
	assign w_sys_tmp3855 = 32'sh000002e8;
	assign w_sys_tmp3860 = (w_sys_tmp3861 + r_run_k_29);
	assign w_sys_tmp3861 = 32'sh00000307;
	assign w_sys_tmp3866 = (w_sys_tmp3867 + r_run_k_29);
	assign w_sys_tmp3867 = 32'sh00000326;
	assign w_sys_tmp3884 = (w_sys_tmp3885 + r_run_k_29);
	assign w_sys_tmp3885 = 32'sh00000345;
	assign w_sys_tmp3890 = (w_sys_tmp3891 + r_run_k_29);
	assign w_sys_tmp3891 = 32'sh00000364;
	assign w_sys_tmp3896 = (w_sys_tmp3897 + r_run_k_29);
	assign w_sys_tmp3897 = 32'sh00000383;
	assign w_sys_tmp3902 = (w_sys_tmp3903 + r_run_k_29);
	assign w_sys_tmp3903 = 32'sh000003a2;
	assign w_sys_tmp3908 = (w_sys_tmp3909 + r_run_k_29);
	assign w_sys_tmp3909 = 32'sh000003c1;
	assign w_sys_tmp3913 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp3914 = 32'sh00000002;
	assign w_sys_tmp3915 = ( !w_sys_tmp3916 );
	assign w_sys_tmp3916 = (w_sys_tmp3917 < r_run_k_29);
	assign w_sys_tmp3917 = 32'sh00000007;
	assign w_sys_tmp3920 = (w_sys_tmp3921 + r_run_k_29);
	assign w_sys_tmp3921 = 32'sh0000003e;
	assign w_sys_tmp3922 = w_sub00_result_dataout;
	assign w_sys_tmp3926 = (w_sys_tmp3927 + r_run_k_29);
	assign w_sys_tmp3927 = 32'sh0000005d;
	assign w_sys_tmp3932 = (w_sys_tmp3933 + r_run_k_29);
	assign w_sys_tmp3933 = 32'sh0000007c;
	assign w_sys_tmp3938 = (w_sys_tmp3939 + r_run_k_29);
	assign w_sys_tmp3939 = 32'sh0000009b;
	assign w_sys_tmp3944 = (w_sys_tmp3945 + r_run_k_29);
	assign w_sys_tmp3945 = 32'sh000000ba;
	assign w_sys_tmp3950 = (w_sys_tmp3951 + r_run_k_29);
	assign w_sys_tmp3951 = 32'sh000000d9;
	assign w_sys_tmp3956 = (w_sys_tmp3957 + r_run_k_29);
	assign w_sys_tmp3957 = 32'sh000000f8;
	assign w_sys_tmp3961 = (w_sys_tmp3962 + r_run_k_29);
	assign w_sys_tmp3962 = 32'sh00000117;
	assign w_sys_tmp3966 = (w_sys_tmp3967 + r_run_k_29);
	assign w_sys_tmp3967 = 32'sh00000136;
	assign w_sys_tmp3971 = (w_sys_tmp3972 + r_run_k_29);
	assign w_sys_tmp3972 = 32'sh00000155;
	assign w_sys_tmp3976 = (w_sys_tmp3977 + r_run_k_29);
	assign w_sys_tmp3977 = 32'sh00000174;
	assign w_sys_tmp3981 = (w_sys_tmp3982 + r_run_k_29);
	assign w_sys_tmp3982 = 32'sh00000193;
	assign w_sys_tmp3986 = (w_sys_tmp3987 + r_run_k_29);
	assign w_sys_tmp3987 = 32'sh000001b2;
	assign w_sys_tmp3991 = (w_sys_tmp3992 + r_run_k_29);
	assign w_sys_tmp3992 = 32'sh000001d1;
	assign w_sys_tmp3996 = (w_sys_tmp3997 + r_run_k_29);
	assign w_sys_tmp3997 = 32'sh000001f0;
	assign w_sys_tmp4001 = (w_sys_tmp4002 + r_run_k_29);
	assign w_sys_tmp4002 = 32'sh0000020f;
	assign w_sys_tmp4006 = (w_sys_tmp4007 + r_run_k_29);
	assign w_sys_tmp4007 = 32'sh0000022e;
	assign w_sys_tmp4011 = (w_sys_tmp4012 + r_run_k_29);
	assign w_sys_tmp4012 = 32'sh0000024d;
	assign w_sys_tmp4016 = (w_sys_tmp4017 + r_run_k_29);
	assign w_sys_tmp4017 = 32'sh0000026c;
	assign w_sys_tmp4021 = (w_sys_tmp4022 + r_run_k_29);
	assign w_sys_tmp4022 = 32'sh0000028b;
	assign w_sys_tmp4026 = (w_sys_tmp4027 + r_run_k_29);
	assign w_sys_tmp4027 = 32'sh000002aa;
	assign w_sys_tmp4031 = (w_sys_tmp4032 + r_run_k_29);
	assign w_sys_tmp4032 = 32'sh000002c9;
	assign w_sys_tmp4036 = (w_sys_tmp4037 + r_run_k_29);
	assign w_sys_tmp4037 = 32'sh000002e8;
	assign w_sys_tmp4041 = (w_sys_tmp4042 + r_run_k_29);
	assign w_sys_tmp4042 = 32'sh00000307;
	assign w_sys_tmp4046 = (w_sys_tmp4047 + r_run_k_29);
	assign w_sys_tmp4047 = 32'sh00000326;
	assign w_sys_tmp4051 = (w_sys_tmp4052 + r_run_k_29);
	assign w_sys_tmp4052 = 32'sh00000345;
	assign w_sys_tmp4056 = (w_sys_tmp4057 + r_run_k_29);
	assign w_sys_tmp4057 = 32'sh00000364;
	assign w_sys_tmp4061 = (w_sys_tmp4062 + r_run_k_29);
	assign w_sys_tmp4062 = 32'sh00000383;
	assign w_sys_tmp4066 = (w_sys_tmp4067 + r_run_k_29);
	assign w_sys_tmp4067 = 32'sh000003a2;
	assign w_sys_tmp4071 = (w_sys_tmp4072 + r_run_k_29);
	assign w_sys_tmp4072 = 32'sh00000044;
	assign w_sys_tmp4076 = (w_sys_tmp4077 + r_run_k_29);
	assign w_sys_tmp4077 = 32'sh00000063;
	assign w_sys_tmp4081 = (w_sys_tmp4082 + r_run_k_29);
	assign w_sys_tmp4082 = 32'sh00000082;
	assign w_sys_tmp4086 = (w_sys_tmp4087 + r_run_k_29);
	assign w_sys_tmp4087 = 32'sh000000a1;
	assign w_sys_tmp4091 = (w_sys_tmp4092 + r_run_k_29);
	assign w_sys_tmp4092 = 32'sh000000c0;
	assign w_sys_tmp4096 = (w_sys_tmp4097 + r_run_k_29);
	assign w_sys_tmp4097 = 32'sh000000df;
	assign w_sys_tmp4101 = (w_sys_tmp4102 + r_run_k_29);
	assign w_sys_tmp4102 = 32'sh000000fe;
	assign w_sys_tmp4106 = (w_sys_tmp4107 + r_run_k_29);
	assign w_sys_tmp4107 = 32'sh0000011d;
	assign w_sys_tmp4111 = (w_sys_tmp4112 + r_run_k_29);
	assign w_sys_tmp4112 = 32'sh0000013c;
	assign w_sys_tmp4116 = (w_sys_tmp4117 + r_run_k_29);
	assign w_sys_tmp4117 = 32'sh0000015b;
	assign w_sys_tmp4121 = (w_sys_tmp4122 + r_run_k_29);
	assign w_sys_tmp4122 = 32'sh0000017a;
	assign w_sys_tmp4126 = (w_sys_tmp4127 + r_run_k_29);
	assign w_sys_tmp4127 = 32'sh00000199;
	assign w_sys_tmp4131 = (w_sys_tmp4132 + r_run_k_29);
	assign w_sys_tmp4132 = 32'sh000001b8;
	assign w_sys_tmp4136 = (w_sys_tmp4137 + r_run_k_29);
	assign w_sys_tmp4137 = 32'sh000001d7;
	assign w_sys_tmp4141 = (w_sys_tmp4142 + r_run_k_29);
	assign w_sys_tmp4142 = 32'sh000001f6;
	assign w_sys_tmp4146 = (w_sys_tmp4147 + r_run_k_29);
	assign w_sys_tmp4147 = 32'sh00000215;
	assign w_sys_tmp4151 = (w_sys_tmp4152 + r_run_k_29);
	assign w_sys_tmp4152 = 32'sh00000234;
	assign w_sys_tmp4156 = (w_sys_tmp4157 + r_run_k_29);
	assign w_sys_tmp4157 = 32'sh00000253;
	assign w_sys_tmp4161 = (w_sys_tmp4162 + r_run_k_29);
	assign w_sys_tmp4162 = 32'sh00000272;
	assign w_sys_tmp4166 = (w_sys_tmp4167 + r_run_k_29);
	assign w_sys_tmp4167 = 32'sh00000291;
	assign w_sys_tmp4171 = (w_sys_tmp4172 + r_run_k_29);
	assign w_sys_tmp4172 = 32'sh000002b0;
	assign w_sys_tmp4176 = (w_sys_tmp4177 + r_run_k_29);
	assign w_sys_tmp4177 = 32'sh000002cf;
	assign w_sys_tmp4181 = (w_sys_tmp4182 + r_run_k_29);
	assign w_sys_tmp4182 = 32'sh000002ee;
	assign w_sys_tmp4186 = (w_sys_tmp4187 + r_run_k_29);
	assign w_sys_tmp4187 = 32'sh0000030d;
	assign w_sys_tmp4191 = (w_sys_tmp4192 + r_run_k_29);
	assign w_sys_tmp4192 = 32'sh0000032c;
	assign w_sys_tmp4196 = (w_sys_tmp4197 + r_run_k_29);
	assign w_sys_tmp4197 = 32'sh0000034b;
	assign w_sys_tmp4201 = (w_sys_tmp4202 + r_run_k_29);
	assign w_sys_tmp4202 = 32'sh0000036a;
	assign w_sys_tmp4206 = (w_sys_tmp4207 + r_run_k_29);
	assign w_sys_tmp4207 = 32'sh00000389;
	assign w_sys_tmp4211 = (w_sys_tmp4212 + r_run_k_29);
	assign w_sys_tmp4212 = 32'sh000003a8;
	assign w_sys_tmp4216 = (w_sys_tmp4217 + r_run_k_29);
	assign w_sys_tmp4217 = 32'sh0000004a;
	assign w_sys_tmp4221 = (w_sys_tmp4222 + r_run_k_29);
	assign w_sys_tmp4222 = 32'sh00000069;
	assign w_sys_tmp4226 = (w_sys_tmp4227 + r_run_k_29);
	assign w_sys_tmp4227 = 32'sh00000088;
	assign w_sys_tmp4231 = (w_sys_tmp4232 + r_run_k_29);
	assign w_sys_tmp4232 = 32'sh000000a7;
	assign w_sys_tmp4236 = (w_sys_tmp4237 + r_run_k_29);
	assign w_sys_tmp4237 = 32'sh000000c6;
	assign w_sys_tmp4241 = (w_sys_tmp4242 + r_run_k_29);
	assign w_sys_tmp4242 = 32'sh000000e5;
	assign w_sys_tmp4246 = (w_sys_tmp4247 + r_run_k_29);
	assign w_sys_tmp4247 = 32'sh00000104;
	assign w_sys_tmp4251 = (w_sys_tmp4252 + r_run_k_29);
	assign w_sys_tmp4252 = 32'sh00000123;
	assign w_sys_tmp4256 = (w_sys_tmp4257 + r_run_k_29);
	assign w_sys_tmp4257 = 32'sh00000142;
	assign w_sys_tmp4261 = (w_sys_tmp4262 + r_run_k_29);
	assign w_sys_tmp4262 = 32'sh00000161;
	assign w_sys_tmp4266 = (w_sys_tmp4267 + r_run_k_29);
	assign w_sys_tmp4267 = 32'sh00000180;
	assign w_sys_tmp4271 = (w_sys_tmp4272 + r_run_k_29);
	assign w_sys_tmp4272 = 32'sh0000019f;
	assign w_sys_tmp4276 = (w_sys_tmp4277 + r_run_k_29);
	assign w_sys_tmp4277 = 32'sh000001be;
	assign w_sys_tmp4281 = (w_sys_tmp4282 + r_run_k_29);
	assign w_sys_tmp4282 = 32'sh000001dd;
	assign w_sys_tmp4286 = (w_sys_tmp4287 + r_run_k_29);
	assign w_sys_tmp4287 = 32'sh000001fc;
	assign w_sys_tmp4291 = (w_sys_tmp4292 + r_run_k_29);
	assign w_sys_tmp4292 = 32'sh0000021b;
	assign w_sys_tmp4296 = (w_sys_tmp4297 + r_run_k_29);
	assign w_sys_tmp4297 = 32'sh0000023a;
	assign w_sys_tmp4301 = (w_sys_tmp4302 + r_run_k_29);
	assign w_sys_tmp4302 = 32'sh00000259;
	assign w_sys_tmp4306 = (w_sys_tmp4307 + r_run_k_29);
	assign w_sys_tmp4307 = 32'sh00000278;
	assign w_sys_tmp4311 = (w_sys_tmp4312 + r_run_k_29);
	assign w_sys_tmp4312 = 32'sh00000297;
	assign w_sys_tmp4316 = (w_sys_tmp4317 + r_run_k_29);
	assign w_sys_tmp4317 = 32'sh000002b6;
	assign w_sys_tmp4321 = (w_sys_tmp4322 + r_run_k_29);
	assign w_sys_tmp4322 = 32'sh000002d5;
	assign w_sys_tmp4326 = (w_sys_tmp4327 + r_run_k_29);
	assign w_sys_tmp4327 = 32'sh000002f4;
	assign w_sys_tmp4331 = (w_sys_tmp4332 + r_run_k_29);
	assign w_sys_tmp4332 = 32'sh00000313;
	assign w_sys_tmp4336 = (w_sys_tmp4337 + r_run_k_29);
	assign w_sys_tmp4337 = 32'sh00000332;
	assign w_sys_tmp4341 = (w_sys_tmp4342 + r_run_k_29);
	assign w_sys_tmp4342 = 32'sh00000351;
	assign w_sys_tmp4346 = (w_sys_tmp4347 + r_run_k_29);
	assign w_sys_tmp4347 = 32'sh00000370;
	assign w_sys_tmp4351 = (w_sys_tmp4352 + r_run_k_29);
	assign w_sys_tmp4352 = 32'sh0000038f;
	assign w_sys_tmp4356 = (w_sys_tmp4357 + r_run_k_29);
	assign w_sys_tmp4357 = 32'sh000003ae;
	assign w_sys_tmp4361 = (w_sys_tmp4362 + r_run_k_29);
	assign w_sys_tmp4362 = 32'sh00000050;
	assign w_sys_tmp4366 = (w_sys_tmp4367 + r_run_k_29);
	assign w_sys_tmp4367 = 32'sh0000006f;
	assign w_sys_tmp4371 = (w_sys_tmp4372 + r_run_k_29);
	assign w_sys_tmp4372 = 32'sh0000008e;
	assign w_sys_tmp4376 = (w_sys_tmp4377 + r_run_k_29);
	assign w_sys_tmp4377 = 32'sh000000ad;
	assign w_sys_tmp4381 = (w_sys_tmp4382 + r_run_k_29);
	assign w_sys_tmp4382 = 32'sh000000cc;
	assign w_sys_tmp4386 = (w_sys_tmp4387 + r_run_k_29);
	assign w_sys_tmp4387 = 32'sh000000eb;
	assign w_sys_tmp4391 = (w_sys_tmp4392 + r_run_k_29);
	assign w_sys_tmp4392 = 32'sh0000010a;
	assign w_sys_tmp4396 = (w_sys_tmp4397 + r_run_k_29);
	assign w_sys_tmp4397 = 32'sh00000129;
	assign w_sys_tmp4401 = (w_sys_tmp4402 + r_run_k_29);
	assign w_sys_tmp4402 = 32'sh00000148;
	assign w_sys_tmp4406 = (w_sys_tmp4407 + r_run_k_29);
	assign w_sys_tmp4407 = 32'sh00000167;
	assign w_sys_tmp4411 = (w_sys_tmp4412 + r_run_k_29);
	assign w_sys_tmp4412 = 32'sh00000186;
	assign w_sys_tmp4416 = (w_sys_tmp4417 + r_run_k_29);
	assign w_sys_tmp4417 = 32'sh000001a5;
	assign w_sys_tmp4421 = (w_sys_tmp4422 + r_run_k_29);
	assign w_sys_tmp4422 = 32'sh000001c4;
	assign w_sys_tmp4426 = (w_sys_tmp4427 + r_run_k_29);
	assign w_sys_tmp4427 = 32'sh000001e3;
	assign w_sys_tmp4431 = (w_sys_tmp4432 + r_run_k_29);
	assign w_sys_tmp4432 = 32'sh00000202;
	assign w_sys_tmp4436 = (w_sys_tmp4437 + r_run_k_29);
	assign w_sys_tmp4437 = 32'sh00000221;
	assign w_sys_tmp4441 = (w_sys_tmp4442 + r_run_k_29);
	assign w_sys_tmp4442 = 32'sh00000240;
	assign w_sys_tmp4446 = (w_sys_tmp4447 + r_run_k_29);
	assign w_sys_tmp4447 = 32'sh0000025f;
	assign w_sys_tmp4451 = (w_sys_tmp4452 + r_run_k_29);
	assign w_sys_tmp4452 = 32'sh0000027e;
	assign w_sys_tmp4456 = (w_sys_tmp4457 + r_run_k_29);
	assign w_sys_tmp4457 = 32'sh0000029d;
	assign w_sys_tmp4461 = (w_sys_tmp4462 + r_run_k_29);
	assign w_sys_tmp4462 = 32'sh000002bc;
	assign w_sys_tmp4466 = (w_sys_tmp4467 + r_run_k_29);
	assign w_sys_tmp4467 = 32'sh000002db;
	assign w_sys_tmp4471 = (w_sys_tmp4472 + r_run_k_29);
	assign w_sys_tmp4472 = 32'sh000002fa;
	assign w_sys_tmp4476 = (w_sys_tmp4477 + r_run_k_29);
	assign w_sys_tmp4477 = 32'sh00000319;
	assign w_sys_tmp4481 = (w_sys_tmp4482 + r_run_k_29);
	assign w_sys_tmp4482 = 32'sh00000338;
	assign w_sys_tmp4486 = (w_sys_tmp4487 + r_run_k_29);
	assign w_sys_tmp4487 = 32'sh00000357;
	assign w_sys_tmp4491 = (w_sys_tmp4492 + r_run_k_29);
	assign w_sys_tmp4492 = 32'sh00000376;
	assign w_sys_tmp4496 = (w_sys_tmp4497 + r_run_k_29);
	assign w_sys_tmp4497 = 32'sh00000395;
	assign w_sys_tmp4501 = (w_sys_tmp4502 + r_run_k_29);
	assign w_sys_tmp4502 = 32'sh000003b4;
	assign w_sys_tmp4505 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp4506 = 32'sh0000001a;
	assign w_sys_tmp4507 = ( !w_sys_tmp4508 );
	assign w_sys_tmp4508 = (w_sys_tmp4509 < r_run_k_29);
	assign w_sys_tmp4509 = 32'sh0000001e;
	assign w_sys_tmp4512 = (w_sys_tmp4513 + r_run_k_29);
	assign w_sys_tmp4513 = 32'sh0000003e;
	assign w_sys_tmp4514 = w_sub20_result_dataout;
	assign w_sys_tmp4518 = (w_sys_tmp4519 + r_run_k_29);
	assign w_sys_tmp4519 = 32'sh0000005d;
	assign w_sys_tmp4524 = (w_sys_tmp4525 + r_run_k_29);
	assign w_sys_tmp4525 = 32'sh0000007c;
	assign w_sys_tmp4530 = (w_sys_tmp4531 + r_run_k_29);
	assign w_sys_tmp4531 = 32'sh0000009b;
	assign w_sys_tmp4536 = (w_sys_tmp4537 + r_run_k_29);
	assign w_sys_tmp4537 = 32'sh000000ba;
	assign w_sys_tmp4542 = (w_sys_tmp4543 + r_run_k_29);
	assign w_sys_tmp4543 = 32'sh000000d9;
	assign w_sys_tmp4548 = (w_sys_tmp4549 + r_run_k_29);
	assign w_sys_tmp4549 = 32'sh000000f8;
	assign w_sys_tmp4553 = (w_sys_tmp4554 + r_run_k_29);
	assign w_sys_tmp4554 = 32'sh00000117;
	assign w_sys_tmp4558 = (w_sys_tmp4559 + r_run_k_29);
	assign w_sys_tmp4559 = 32'sh00000136;
	assign w_sys_tmp4563 = (w_sys_tmp4564 + r_run_k_29);
	assign w_sys_tmp4564 = 32'sh00000155;
	assign w_sys_tmp4568 = (w_sys_tmp4569 + r_run_k_29);
	assign w_sys_tmp4569 = 32'sh00000174;
	assign w_sys_tmp4573 = (w_sys_tmp4574 + r_run_k_29);
	assign w_sys_tmp4574 = 32'sh00000193;
	assign w_sys_tmp4578 = (w_sys_tmp4579 + r_run_k_29);
	assign w_sys_tmp4579 = 32'sh000001b2;
	assign w_sys_tmp4583 = (w_sys_tmp4584 + r_run_k_29);
	assign w_sys_tmp4584 = 32'sh000001d1;
	assign w_sys_tmp4588 = (w_sys_tmp4589 + r_run_k_29);
	assign w_sys_tmp4589 = 32'sh000001f0;
	assign w_sys_tmp4593 = (w_sys_tmp4594 + r_run_k_29);
	assign w_sys_tmp4594 = 32'sh0000020f;
	assign w_sys_tmp4598 = (w_sys_tmp4599 + r_run_k_29);
	assign w_sys_tmp4599 = 32'sh0000022e;
	assign w_sys_tmp4603 = (w_sys_tmp4604 + r_run_k_29);
	assign w_sys_tmp4604 = 32'sh0000024d;
	assign w_sys_tmp4608 = (w_sys_tmp4609 + r_run_k_29);
	assign w_sys_tmp4609 = 32'sh0000026c;
	assign w_sys_tmp4613 = (w_sys_tmp4614 + r_run_k_29);
	assign w_sys_tmp4614 = 32'sh0000028b;
	assign w_sys_tmp4618 = (w_sys_tmp4619 + r_run_k_29);
	assign w_sys_tmp4619 = 32'sh000002aa;
	assign w_sys_tmp4623 = (w_sys_tmp4624 + r_run_k_29);
	assign w_sys_tmp4624 = 32'sh000002c9;
	assign w_sys_tmp4628 = (w_sys_tmp4629 + r_run_k_29);
	assign w_sys_tmp4629 = 32'sh000002e8;
	assign w_sys_tmp4633 = (w_sys_tmp4634 + r_run_k_29);
	assign w_sys_tmp4634 = 32'sh00000307;
	assign w_sys_tmp4638 = (w_sys_tmp4639 + r_run_k_29);
	assign w_sys_tmp4639 = 32'sh00000326;
	assign w_sys_tmp4643 = (w_sys_tmp4644 + r_run_k_29);
	assign w_sys_tmp4644 = 32'sh00000345;
	assign w_sys_tmp4648 = (w_sys_tmp4649 + r_run_k_29);
	assign w_sys_tmp4649 = 32'sh00000364;
	assign w_sys_tmp4653 = (w_sys_tmp4654 + r_run_k_29);
	assign w_sys_tmp4654 = 32'sh00000383;
	assign w_sys_tmp4658 = (w_sys_tmp4659 + r_run_k_29);
	assign w_sys_tmp4659 = 32'sh000003a2;
	assign w_sys_tmp4662 = (r_run_k_29 + w_sys_intOne);


	sub19
		sub19_inst(
			.i_fld_T_0_addr_0 (w_sub19_T_addr),
			.i_fld_T_0_datain_0 (w_sub19_T_datain),
			.o_fld_T_0_dataout_0 (w_sub19_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub19_T_r_w),
			.i_fld_U_2_addr_0 (w_sub19_U_addr),
			.i_fld_U_2_datain_0 (w_sub19_U_datain),
			.o_fld_U_2_dataout_0 (w_sub19_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub19_U_r_w),
			.i_fld_V_1_addr_0 (w_sub19_V_addr),
			.i_fld_V_1_datain_0 (w_sub19_V_datain),
			.o_fld_V_1_dataout_0 (w_sub19_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub19_V_r_w),
			.i_fld_result_3_addr_0 (w_sub19_result_addr),
			.i_fld_result_3_datain_0 (w_sub19_result_datain),
			.o_fld_result_3_dataout_0 (w_sub19_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub19_result_r_w),
			.o_run_busy (w_sub19_run_busy),
			.i_run_req (r_sub19_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub09
		sub09_inst(
			.i_fld_T_0_addr_0 (w_sub09_T_addr),
			.i_fld_T_0_datain_0 (w_sub09_T_datain),
			.o_fld_T_0_dataout_0 (w_sub09_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub09_T_r_w),
			.i_fld_U_2_addr_0 (w_sub09_U_addr),
			.i_fld_U_2_datain_0 (w_sub09_U_datain),
			.o_fld_U_2_dataout_0 (w_sub09_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub09_U_r_w),
			.i_fld_V_1_addr_0 (w_sub09_V_addr),
			.i_fld_V_1_datain_0 (w_sub09_V_datain),
			.o_fld_V_1_dataout_0 (w_sub09_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub09_V_r_w),
			.i_fld_result_3_addr_0 (w_sub09_result_addr),
			.i_fld_result_3_datain_0 (w_sub09_result_datain),
			.o_fld_result_3_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub09_result_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_T_0_addr_0 (w_sub08_T_addr),
			.i_fld_T_0_datain_0 (w_sub08_T_datain),
			.o_fld_T_0_dataout_0 (w_sub08_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub08_T_r_w),
			.i_fld_U_2_addr_0 (w_sub08_U_addr),
			.i_fld_U_2_datain_0 (w_sub08_U_datain),
			.o_fld_U_2_dataout_0 (w_sub08_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub08_U_r_w),
			.i_fld_V_1_addr_0 (w_sub08_V_addr),
			.i_fld_V_1_datain_0 (w_sub08_V_datain),
			.o_fld_V_1_dataout_0 (w_sub08_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub08_V_r_w),
			.i_fld_result_3_addr_0 (w_sub08_result_addr),
			.i_fld_result_3_datain_0 (w_sub08_result_datain),
			.o_fld_result_3_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub08_result_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub24
		sub24_inst(
			.i_fld_T_0_addr_0 (w_sub24_T_addr),
			.i_fld_T_0_datain_0 (w_sub24_T_datain),
			.o_fld_T_0_dataout_0 (w_sub24_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub24_T_r_w),
			.i_fld_U_2_addr_0 (w_sub24_U_addr),
			.i_fld_U_2_datain_0 (w_sub24_U_datain),
			.o_fld_U_2_dataout_0 (w_sub24_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub24_U_r_w),
			.i_fld_V_1_addr_0 (w_sub24_V_addr),
			.i_fld_V_1_datain_0 (w_sub24_V_datain),
			.o_fld_V_1_dataout_0 (w_sub24_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub24_V_r_w),
			.i_fld_result_3_addr_0 (w_sub24_result_addr),
			.i_fld_result_3_datain_0 (w_sub24_result_datain),
			.o_fld_result_3_dataout_0 (w_sub24_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub24_result_r_w),
			.o_run_busy (w_sub24_run_busy),
			.i_run_req (r_sub24_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub22
		sub22_inst(
			.i_fld_T_0_addr_0 (w_sub22_T_addr),
			.i_fld_T_0_datain_0 (w_sub22_T_datain),
			.o_fld_T_0_dataout_0 (w_sub22_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub22_T_r_w),
			.i_fld_U_2_addr_0 (w_sub22_U_addr),
			.i_fld_U_2_datain_0 (w_sub22_U_datain),
			.o_fld_U_2_dataout_0 (w_sub22_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub22_U_r_w),
			.i_fld_V_1_addr_0 (w_sub22_V_addr),
			.i_fld_V_1_datain_0 (w_sub22_V_datain),
			.o_fld_V_1_dataout_0 (w_sub22_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub22_V_r_w),
			.i_fld_result_3_addr_0 (w_sub22_result_addr),
			.i_fld_result_3_datain_0 (w_sub22_result_datain),
			.o_fld_result_3_dataout_0 (w_sub22_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub22_result_r_w),
			.o_run_busy (w_sub22_run_busy),
			.i_run_req (r_sub22_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub23
		sub23_inst(
			.i_fld_T_0_addr_0 (w_sub23_T_addr),
			.i_fld_T_0_datain_0 (w_sub23_T_datain),
			.o_fld_T_0_dataout_0 (w_sub23_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub23_T_r_w),
			.i_fld_U_2_addr_0 (w_sub23_U_addr),
			.i_fld_U_2_datain_0 (w_sub23_U_datain),
			.o_fld_U_2_dataout_0 (w_sub23_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub23_U_r_w),
			.i_fld_V_1_addr_0 (w_sub23_V_addr),
			.i_fld_V_1_datain_0 (w_sub23_V_datain),
			.o_fld_V_1_dataout_0 (w_sub23_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub23_V_r_w),
			.i_fld_result_3_addr_0 (w_sub23_result_addr),
			.i_fld_result_3_datain_0 (w_sub23_result_datain),
			.o_fld_result_3_dataout_0 (w_sub23_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub23_result_r_w),
			.o_run_busy (w_sub23_run_busy),
			.i_run_req (r_sub23_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_T_0_addr_0 (w_sub12_T_addr),
			.i_fld_T_0_datain_0 (w_sub12_T_datain),
			.o_fld_T_0_dataout_0 (w_sub12_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub12_T_r_w),
			.i_fld_U_2_addr_0 (w_sub12_U_addr),
			.i_fld_U_2_datain_0 (w_sub12_U_datain),
			.o_fld_U_2_dataout_0 (w_sub12_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub12_U_r_w),
			.i_fld_V_1_addr_0 (w_sub12_V_addr),
			.i_fld_V_1_datain_0 (w_sub12_V_datain),
			.o_fld_V_1_dataout_0 (w_sub12_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub12_V_r_w),
			.i_fld_result_3_addr_0 (w_sub12_result_addr),
			.i_fld_result_3_datain_0 (w_sub12_result_datain),
			.o_fld_result_3_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub12_result_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_T_0_addr_0 (w_sub03_T_addr),
			.i_fld_T_0_datain_0 (w_sub03_T_datain),
			.o_fld_T_0_dataout_0 (w_sub03_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub03_T_r_w),
			.i_fld_U_2_addr_0 (w_sub03_U_addr),
			.i_fld_U_2_datain_0 (w_sub03_U_datain),
			.o_fld_U_2_dataout_0 (w_sub03_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub03_U_r_w),
			.i_fld_V_1_addr_0 (w_sub03_V_addr),
			.i_fld_V_1_datain_0 (w_sub03_V_datain),
			.o_fld_V_1_dataout_0 (w_sub03_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub03_V_r_w),
			.i_fld_result_3_addr_0 (w_sub03_result_addr),
			.i_fld_result_3_datain_0 (w_sub03_result_datain),
			.o_fld_result_3_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub03_result_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_T_0_addr_0 (w_sub02_T_addr),
			.i_fld_T_0_datain_0 (w_sub02_T_datain),
			.o_fld_T_0_dataout_0 (w_sub02_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub02_T_r_w),
			.i_fld_U_2_addr_0 (w_sub02_U_addr),
			.i_fld_U_2_datain_0 (w_sub02_U_datain),
			.o_fld_U_2_dataout_0 (w_sub02_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub02_U_r_w),
			.i_fld_V_1_addr_0 (w_sub02_V_addr),
			.i_fld_V_1_datain_0 (w_sub02_V_datain),
			.o_fld_V_1_dataout_0 (w_sub02_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub02_V_r_w),
			.i_fld_result_3_addr_0 (w_sub02_result_addr),
			.i_fld_result_3_datain_0 (w_sub02_result_datain),
			.o_fld_result_3_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub02_result_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_T_0_addr_0 (w_sub11_T_addr),
			.i_fld_T_0_datain_0 (w_sub11_T_datain),
			.o_fld_T_0_dataout_0 (w_sub11_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub11_T_r_w),
			.i_fld_U_2_addr_0 (w_sub11_U_addr),
			.i_fld_U_2_datain_0 (w_sub11_U_datain),
			.o_fld_U_2_dataout_0 (w_sub11_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub11_U_r_w),
			.i_fld_V_1_addr_0 (w_sub11_V_addr),
			.i_fld_V_1_datain_0 (w_sub11_V_datain),
			.o_fld_V_1_dataout_0 (w_sub11_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub11_V_r_w),
			.i_fld_result_3_addr_0 (w_sub11_result_addr),
			.i_fld_result_3_datain_0 (w_sub11_result_datain),
			.o_fld_result_3_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub11_result_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_T_0_addr_0 (w_sub14_T_addr),
			.i_fld_T_0_datain_0 (w_sub14_T_datain),
			.o_fld_T_0_dataout_0 (w_sub14_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub14_T_r_w),
			.i_fld_U_2_addr_0 (w_sub14_U_addr),
			.i_fld_U_2_datain_0 (w_sub14_U_datain),
			.o_fld_U_2_dataout_0 (w_sub14_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub14_U_r_w),
			.i_fld_V_1_addr_0 (w_sub14_V_addr),
			.i_fld_V_1_datain_0 (w_sub14_V_datain),
			.o_fld_V_1_dataout_0 (w_sub14_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub14_V_r_w),
			.i_fld_result_3_addr_0 (w_sub14_result_addr),
			.i_fld_result_3_datain_0 (w_sub14_result_datain),
			.o_fld_result_3_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub14_result_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_T_0_addr_0 (w_sub01_T_addr),
			.i_fld_T_0_datain_0 (w_sub01_T_datain),
			.o_fld_T_0_dataout_0 (w_sub01_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub01_T_r_w),
			.i_fld_U_2_addr_0 (w_sub01_U_addr),
			.i_fld_U_2_datain_0 (w_sub01_U_datain),
			.o_fld_U_2_dataout_0 (w_sub01_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub01_U_r_w),
			.i_fld_V_1_addr_0 (w_sub01_V_addr),
			.i_fld_V_1_datain_0 (w_sub01_V_datain),
			.o_fld_V_1_dataout_0 (w_sub01_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub01_V_r_w),
			.i_fld_result_3_addr_0 (w_sub01_result_addr),
			.i_fld_result_3_datain_0 (w_sub01_result_datain),
			.o_fld_result_3_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub01_result_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_T_0_addr_0 (w_sub00_T_addr),
			.i_fld_T_0_datain_0 (w_sub00_T_datain),
			.o_fld_T_0_dataout_0 (w_sub00_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub00_T_r_w),
			.i_fld_U_2_addr_0 (w_sub00_U_addr),
			.i_fld_U_2_datain_0 (w_sub00_U_datain),
			.o_fld_U_2_dataout_0 (w_sub00_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub00_U_r_w),
			.i_fld_V_1_addr_0 (w_sub00_V_addr),
			.i_fld_V_1_datain_0 (w_sub00_V_datain),
			.o_fld_V_1_dataout_0 (w_sub00_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub00_V_r_w),
			.i_fld_result_3_addr_0 (w_sub00_result_addr),
			.i_fld_result_3_datain_0 (w_sub00_result_datain),
			.o_fld_result_3_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub00_result_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_T_0_addr_0 (w_sub13_T_addr),
			.i_fld_T_0_datain_0 (w_sub13_T_datain),
			.o_fld_T_0_dataout_0 (w_sub13_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub13_T_r_w),
			.i_fld_U_2_addr_0 (w_sub13_U_addr),
			.i_fld_U_2_datain_0 (w_sub13_U_datain),
			.o_fld_U_2_dataout_0 (w_sub13_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub13_U_r_w),
			.i_fld_V_1_addr_0 (w_sub13_V_addr),
			.i_fld_V_1_datain_0 (w_sub13_V_datain),
			.o_fld_V_1_dataout_0 (w_sub13_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub13_V_r_w),
			.i_fld_result_3_addr_0 (w_sub13_result_addr),
			.i_fld_result_3_datain_0 (w_sub13_result_datain),
			.o_fld_result_3_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub13_result_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_T_0_addr_0 (w_sub07_T_addr),
			.i_fld_T_0_datain_0 (w_sub07_T_datain),
			.o_fld_T_0_dataout_0 (w_sub07_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub07_T_r_w),
			.i_fld_U_2_addr_0 (w_sub07_U_addr),
			.i_fld_U_2_datain_0 (w_sub07_U_datain),
			.o_fld_U_2_dataout_0 (w_sub07_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub07_U_r_w),
			.i_fld_V_1_addr_0 (w_sub07_V_addr),
			.i_fld_V_1_datain_0 (w_sub07_V_datain),
			.o_fld_V_1_dataout_0 (w_sub07_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub07_V_r_w),
			.i_fld_result_3_addr_0 (w_sub07_result_addr),
			.i_fld_result_3_datain_0 (w_sub07_result_datain),
			.o_fld_result_3_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub07_result_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub16
		sub16_inst(
			.i_fld_T_0_addr_0 (w_sub16_T_addr),
			.i_fld_T_0_datain_0 (w_sub16_T_datain),
			.o_fld_T_0_dataout_0 (w_sub16_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub16_T_r_w),
			.i_fld_U_2_addr_0 (w_sub16_U_addr),
			.i_fld_U_2_datain_0 (w_sub16_U_datain),
			.o_fld_U_2_dataout_0 (w_sub16_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub16_U_r_w),
			.i_fld_V_1_addr_0 (w_sub16_V_addr),
			.i_fld_V_1_datain_0 (w_sub16_V_datain),
			.o_fld_V_1_dataout_0 (w_sub16_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub16_V_r_w),
			.i_fld_result_3_addr_0 (w_sub16_result_addr),
			.i_fld_result_3_datain_0 (w_sub16_result_datain),
			.o_fld_result_3_dataout_0 (w_sub16_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub16_result_r_w),
			.o_run_busy (w_sub16_run_busy),
			.i_run_req (r_sub16_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_T_0_addr_0 (w_sub06_T_addr),
			.i_fld_T_0_datain_0 (w_sub06_T_datain),
			.o_fld_T_0_dataout_0 (w_sub06_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub06_T_r_w),
			.i_fld_U_2_addr_0 (w_sub06_U_addr),
			.i_fld_U_2_datain_0 (w_sub06_U_datain),
			.o_fld_U_2_dataout_0 (w_sub06_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub06_U_r_w),
			.i_fld_V_1_addr_0 (w_sub06_V_addr),
			.i_fld_V_1_datain_0 (w_sub06_V_datain),
			.o_fld_V_1_dataout_0 (w_sub06_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub06_V_r_w),
			.i_fld_result_3_addr_0 (w_sub06_result_addr),
			.i_fld_result_3_datain_0 (w_sub06_result_datain),
			.o_fld_result_3_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub06_result_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_T_0_addr_0 (w_sub15_T_addr),
			.i_fld_T_0_datain_0 (w_sub15_T_datain),
			.o_fld_T_0_dataout_0 (w_sub15_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub15_T_r_w),
			.i_fld_U_2_addr_0 (w_sub15_U_addr),
			.i_fld_U_2_datain_0 (w_sub15_U_datain),
			.o_fld_U_2_dataout_0 (w_sub15_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub15_U_r_w),
			.i_fld_V_1_addr_0 (w_sub15_V_addr),
			.i_fld_V_1_datain_0 (w_sub15_V_datain),
			.o_fld_V_1_dataout_0 (w_sub15_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub15_V_r_w),
			.i_fld_result_3_addr_0 (w_sub15_result_addr),
			.i_fld_result_3_datain_0 (w_sub15_result_datain),
			.o_fld_result_3_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub15_result_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_T_0_addr_0 (w_sub05_T_addr),
			.i_fld_T_0_datain_0 (w_sub05_T_datain),
			.o_fld_T_0_dataout_0 (w_sub05_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub05_T_r_w),
			.i_fld_U_2_addr_0 (w_sub05_U_addr),
			.i_fld_U_2_datain_0 (w_sub05_U_datain),
			.o_fld_U_2_dataout_0 (w_sub05_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub05_U_r_w),
			.i_fld_V_1_addr_0 (w_sub05_V_addr),
			.i_fld_V_1_datain_0 (w_sub05_V_datain),
			.o_fld_V_1_dataout_0 (w_sub05_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub05_V_r_w),
			.i_fld_result_3_addr_0 (w_sub05_result_addr),
			.i_fld_result_3_datain_0 (w_sub05_result_datain),
			.o_fld_result_3_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub05_result_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub18
		sub18_inst(
			.i_fld_T_0_addr_0 (w_sub18_T_addr),
			.i_fld_T_0_datain_0 (w_sub18_T_datain),
			.o_fld_T_0_dataout_0 (w_sub18_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub18_T_r_w),
			.i_fld_U_2_addr_0 (w_sub18_U_addr),
			.i_fld_U_2_datain_0 (w_sub18_U_datain),
			.o_fld_U_2_dataout_0 (w_sub18_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub18_U_r_w),
			.i_fld_V_1_addr_0 (w_sub18_V_addr),
			.i_fld_V_1_datain_0 (w_sub18_V_datain),
			.o_fld_V_1_dataout_0 (w_sub18_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub18_V_r_w),
			.i_fld_result_3_addr_0 (w_sub18_result_addr),
			.i_fld_result_3_datain_0 (w_sub18_result_datain),
			.o_fld_result_3_dataout_0 (w_sub18_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub18_result_r_w),
			.o_run_busy (w_sub18_run_busy),
			.i_run_req (r_sub18_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_T_0_addr_0 (w_sub04_T_addr),
			.i_fld_T_0_datain_0 (w_sub04_T_datain),
			.o_fld_T_0_dataout_0 (w_sub04_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub04_T_r_w),
			.i_fld_U_2_addr_0 (w_sub04_U_addr),
			.i_fld_U_2_datain_0 (w_sub04_U_datain),
			.o_fld_U_2_dataout_0 (w_sub04_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub04_U_r_w),
			.i_fld_V_1_addr_0 (w_sub04_V_addr),
			.i_fld_V_1_datain_0 (w_sub04_V_datain),
			.o_fld_V_1_dataout_0 (w_sub04_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub04_V_r_w),
			.i_fld_result_3_addr_0 (w_sub04_result_addr),
			.i_fld_result_3_datain_0 (w_sub04_result_datain),
			.o_fld_result_3_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub04_result_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub17
		sub17_inst(
			.i_fld_T_0_addr_0 (w_sub17_T_addr),
			.i_fld_T_0_datain_0 (w_sub17_T_datain),
			.o_fld_T_0_dataout_0 (w_sub17_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub17_T_r_w),
			.i_fld_U_2_addr_0 (w_sub17_U_addr),
			.i_fld_U_2_datain_0 (w_sub17_U_datain),
			.o_fld_U_2_dataout_0 (w_sub17_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub17_U_r_w),
			.i_fld_V_1_addr_0 (w_sub17_V_addr),
			.i_fld_V_1_datain_0 (w_sub17_V_datain),
			.o_fld_V_1_dataout_0 (w_sub17_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub17_V_r_w),
			.i_fld_result_3_addr_0 (w_sub17_result_addr),
			.i_fld_result_3_datain_0 (w_sub17_result_datain),
			.o_fld_result_3_dataout_0 (w_sub17_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub17_result_r_w),
			.o_run_busy (w_sub17_run_busy),
			.i_run_req (r_sub17_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_T_0_addr_0 (w_sub10_T_addr),
			.i_fld_T_0_datain_0 (w_sub10_T_datain),
			.o_fld_T_0_dataout_0 (w_sub10_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub10_T_r_w),
			.i_fld_U_2_addr_0 (w_sub10_U_addr),
			.i_fld_U_2_datain_0 (w_sub10_U_datain),
			.o_fld_U_2_dataout_0 (w_sub10_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub10_U_r_w),
			.i_fld_V_1_addr_0 (w_sub10_V_addr),
			.i_fld_V_1_datain_0 (w_sub10_V_datain),
			.o_fld_V_1_dataout_0 (w_sub10_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub10_V_r_w),
			.i_fld_result_3_addr_0 (w_sub10_result_addr),
			.i_fld_result_3_datain_0 (w_sub10_result_datain),
			.o_fld_result_3_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub10_result_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub20
		sub20_inst(
			.i_fld_T_0_addr_0 (w_sub20_T_addr),
			.i_fld_T_0_datain_0 (w_sub20_T_datain),
			.o_fld_T_0_dataout_0 (w_sub20_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub20_T_r_w),
			.i_fld_U_2_addr_0 (w_sub20_U_addr),
			.i_fld_U_2_datain_0 (w_sub20_U_datain),
			.o_fld_U_2_dataout_0 (w_sub20_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub20_U_r_w),
			.i_fld_V_1_addr_0 (w_sub20_V_addr),
			.i_fld_V_1_datain_0 (w_sub20_V_datain),
			.o_fld_V_1_dataout_0 (w_sub20_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub20_V_r_w),
			.i_fld_result_3_addr_0 (w_sub20_result_addr),
			.i_fld_result_3_datain_0 (w_sub20_result_datain),
			.o_fld_result_3_dataout_0 (w_sub20_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub20_result_r_w),
			.o_run_busy (w_sub20_run_busy),
			.i_run_req (r_sub20_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub21
		sub21_inst(
			.i_fld_T_0_addr_0 (w_sub21_T_addr),
			.i_fld_T_0_datain_0 (w_sub21_T_datain),
			.o_fld_T_0_dataout_0 (w_sub21_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub21_T_r_w),
			.i_fld_U_2_addr_0 (w_sub21_U_addr),
			.i_fld_U_2_datain_0 (w_sub21_U_datain),
			.o_fld_U_2_dataout_0 (w_sub21_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub21_U_r_w),
			.i_fld_V_1_addr_0 (w_sub21_V_addr),
			.i_fld_V_1_datain_0 (w_sub21_V_datain),
			.o_fld_V_1_dataout_0 (w_sub21_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub21_V_r_w),
			.i_fld_result_3_addr_0 (w_sub21_result_addr),
			.i_fld_result_3_datain_0 (w_sub21_result_datain),
			.o_fld_result_3_dataout_0 (w_sub21_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub21_result_r_w),
			.o_run_busy (w_sub21_run_busy),
			.i_run_req (r_sub21_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_V_3(
			.clk (clock),
			.ce_0 (w_fld_V_3_ce_0),
			.addr_0 (w_fld_V_3_addr_0),
			.datain_0 (w_fld_V_3_datain_0),
			.dataout_0 (w_fld_V_3_dataout_0),
			.r_w_0 (w_fld_V_3_r_w_0),
			.ce_1 (w_fld_V_3_ce_1),
			.addr_1 (r_fld_V_3_addr_1),
			.datain_1 (r_fld_V_3_datain_1),
			.dataout_1 (w_fld_V_3_dataout_1),
			.r_w_1 (r_fld_V_3_r_w_1)
		);

	DivInt
		DivInt_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.dividend (r_ip_DivInt_dividend_0),
			.divisor (r_ip_DivInt_divisor_0),
			.fractional (w_ip_DivInt_fractional_0),
			.quotient (w_ip_DivInt_quotient_0)
		);

	DivInt
		DivInt_inst_1(
			.clk (clock),
			.ce (w_sys_ce),
			.dividend (r_ip_DivInt_dividend_1),
			.divisor (r_ip_DivInt_divisor_1),
			.fractional (w_ip_DivInt_fractional_1),
			.quotient (w_ip_DivInt_quotient_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_dividend_0 <= r_run_mx_32;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_divisor_0 <= w_sys_tmp2685;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_dividend_1 <= r_run_mx_32;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_DivInt_divisor_1 <= w_sys_tmp2689;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp38;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp36;

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp18;

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
									else
									if((8'h7<=r_sys_run_step && r_sys_run_step<=8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_36;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp37;

									end
									else
									if((8'h7<=r_sys_run_step && r_sys_run_step<=8'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==8'hd) || (r_sys_run_step==8'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_41;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp15) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp226) ? 7'h13 : 7'h15);

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2104) ? 7'h19 : 7'h1b);

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2577) ? 7'h20 : 7'h4d);

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2580) ? 7'h24 : 7'h26);

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2597) ? 7'h2a : 7'h2c);

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_phase <= ((w_sys_tmp2686) ? 7'h30 : 7'h32);

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2733) ? 7'h36 : 7'h38);

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3675) ? 7'h3c : 7'h3d);

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_phase <= 7'h3f;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_phase <= 7'h41;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h42;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3915) ? 7'h45 : 7'h47);

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h75)) begin
										r_sys_run_phase <= 7'h42;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 7'h48;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4507) ? 7'h4b : 7'h1d);

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_run_phase <= 7'h48;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h75)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 8'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h27)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1) || (r_sys_run_step==8'h2)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h27)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h75)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h74)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1d)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h4d: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp22[9:0] );

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2588[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2584[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2592[9:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h2) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2601[9:0] );

									end
									else
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2606[9:0] );

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2692[9:0] );

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2738[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2768[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2990[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3212[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3194[9:0] );

									end
									else
									if((r_sys_run_step==8'h35) || (r_sys_run_step==8'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3056[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3518[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3080[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3290[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2966[9:0] );

									end
									else
									if((r_sys_run_step==8'h64) || (r_sys_run_step==8'h66)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3338[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3362[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3440[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3128[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3506[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2774[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2918[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3266[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3380[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3182[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3284[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2762[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3434[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3560[9:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3230[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2954[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2870[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2984[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2798[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e) || (r_sys_run_step==8'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3014[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2780[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d) || (r_sys_run_step==8'h6f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3392[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2996[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2864[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3224[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3608[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2978[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2822[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3092[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2960[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3218[9:0] );

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3644[9:0] );

									end
									else
									if((r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3482[9:0] );

									end
									else
									if((r_sys_run_step==8'h54) || (r_sys_run_step==8'h56)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3242[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3272[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3410[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2972[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3452[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3146[9:0] );

									end
									else
									if((r_sys_run_step==8'h94) || (r_sys_run_step==8'h96)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3626[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2852[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3548[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3236[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3140[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3200[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3662[9:0] );

									end
									else
									if((r_sys_run_step==8'h84) || (r_sys_run_step==8'h86)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3530[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2756[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2858[9:0] );

									end
									else
									if((r_sys_run_step==8'h55) || (r_sys_run_step==8'h57)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3248[9:0] );

									end
									else
									if((r_sys_run_step==8'h83) || (r_sys_run_step==8'h85)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3524[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3428[9:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3512[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3038[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3326[9:0] );

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3650[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3464[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d) || (r_sys_run_step==8'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3008[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2846[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2906[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3098[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2924[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3044[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3602[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2942[9:0] );

									end
									else
									if((r_sys_run_step==8'h45) || (r_sys_run_step==8'h47)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3152[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3296[9:0] );

									end
									else
									if((r_sys_run_step==8'h65) || (r_sys_run_step==8'h67)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3344[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3314[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2804[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3104[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3596[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3134[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3476[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2750[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3176[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2912[9:0] );

									end
									else
									if((r_sys_run_step==8'h36) || (r_sys_run_step==8'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3062[9:0] );

									end
									else
									if((r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3578[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2948[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3320[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3470[9:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3050[9:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3500[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2876[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2816[9:0] );

									end
									else
									if((r_sys_run_step==8'h93) || (r_sys_run_step==8'h95)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3620[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2744[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2894[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3386[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3002[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3422[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3656[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2828[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e) || (r_sys_run_step==8'h40)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3110[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3416[9:0] );

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3566[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3458[9:0] );

									end
									else
									if((r_sys_run_step==8'h46) || (r_sys_run_step==8'h48)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3158[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3614[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3554[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3368[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3086[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3188[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3032[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3668[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3206[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3332[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3446[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3572[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2900[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3374[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2810[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3278[9:0] );

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3722[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3680[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3800[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3866[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3686[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3692[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3704[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3794[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3902[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3740[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3908[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3884[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3746[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3710[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3716[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3758[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3854[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3752[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3698[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3812[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3890[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3764[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3860[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3806[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3848[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3818[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3788[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3836[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3842[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3896[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3770[9:0] );

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4176[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4361[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4001[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4166[9:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4326[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4396[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4441[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4316[9:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4261[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4356[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3932[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4281[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3938[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3981[9:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4151[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4381[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4206[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4461[9:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4466[9:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4426[9:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4271[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4031[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4406[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4071[9:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4181[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4141[9:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4191[9:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4341[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3926[9:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4391[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4211[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4246[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4046[9:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4351[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3961[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4436[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4026[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4496[9:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4196[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4161[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4411[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4091[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3956[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4041[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4011[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4256[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4201[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4311[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4456[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4021[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4111[9:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4346[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4306[9:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4156[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4296[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4401[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4226[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4126[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4331[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4086[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4146[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4366[9:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4416[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4251[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4061[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4101[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4486[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4121[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4036[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4291[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4501[9:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4336[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4016[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4301[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4476[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4286[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4066[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4371[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4376[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3920[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3991[9:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4431[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4131[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4006[9:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4186[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3950[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4446[9:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4276[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4451[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4321[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4116[9:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4236[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3971[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4491[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4096[9:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4471[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4106[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4056[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4216[9:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4231[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4241[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4051[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4076[9:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4266[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4171[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4136[9:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4386[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4081[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3966[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3986[9:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4421[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4221[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4481[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3944[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3996[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3976[9:0] );

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4603[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4643[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4558[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4658[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4563[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4512[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4608[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4628[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4548[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4598[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4553[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4583[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4578[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4536[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4524[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4573[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4530[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4633[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4638[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4613[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4588[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4568[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4542[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4653[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4618[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4518[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4593[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4648[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4623[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2586;

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2591;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'hd)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2604;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2695;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h66)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp85_float;

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp92_float;

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp74_float;

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp90_float;

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp88_float;

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp89_float;

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp77_float;

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp103_float;

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp94_float;

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp97_float;

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp76_float;

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp96_float;

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp84_float;

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp104_float;

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp81_float;

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp109_float;

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp93_float;

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp95_float;

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp102_float;

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp87_float;

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp100_float;

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp75_float;

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp101_float;

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp91_float;

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp105_float;

									end
									else
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h7)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp3922;

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp78_float;

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp82_float;

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp107_float;

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp98_float;

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp83_float;

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp80_float;

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp108_float;

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp99_float;

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp106_float;

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp35_float;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h7)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp4514;

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp16_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h3)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'hd)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9b)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h26)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h75)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h1e)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp27[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (8'h1c<=r_sys_run_step && r_sys_run_step<=8'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp32[9:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h93) || (r_sys_run_step==8'h95)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1995[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d) || (r_sys_run_step==8'h2f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp771[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp507[9:0] );

									end
									else
									if((r_sys_run_step==8'h94) || (r_sys_run_step==8'h96)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2007[9:0] );

									end
									else
									if((r_sys_run_step==8'h84) || (r_sys_run_step==8'h86)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1815[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1131[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp831[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp663[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1983[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1959[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp459[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp591[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp351[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1647[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1767[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp255[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1179[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1407[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1323[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1335[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1635[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1419[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1587[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1899[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e) || (r_sys_run_step==8'h30)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp783[9:0] );

									end
									else
									if((r_sys_run_step==8'h46) || (r_sys_run_step==8'h48)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1071[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1155[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1599[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e) || (r_sys_run_step==8'h40)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp975[9:0] );

									end
									else
									if((r_sys_run_step==8'h83) || (r_sys_run_step==8'h85)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1803[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp447[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1971[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp567[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1035[9:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1755[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1383[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1695[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp495[9:0] );

									end
									else
									if((r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1911[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp711[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp723[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp363[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp603[9:0] );

									end
									else
									if((r_sys_run_step==8'h55) || (r_sys_run_step==8'h57)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1251[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp543[9:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp855[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp699[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1287[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1107[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp819[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1167[9:0] );

									end
									else
									if((r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1719[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1851[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp651[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp483[9:0] );

									end
									else
									if((r_sys_run_step==8'h36) || (r_sys_run_step==8'h38)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp879[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp843[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp675[9:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1215[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp375[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp579[9:0] );

									end
									else
									if((r_sys_run_step==8'h54) || (r_sys_run_step==8'h56)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1239[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1863[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2067[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1611[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp555[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1011[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1659[9:0] );

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2043[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1395[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp639[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1227[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1623[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp735[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1191[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp315[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2091[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp915[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1479[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp231[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1527[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1683[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1143[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp411[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1791[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp243[9:0] );

									end
									else
									if((r_sys_run_step==8'h35) || (r_sys_run_step==8'h37)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp867[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1947[9:0] );

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1887[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1347[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp939[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp927[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d) || (r_sys_run_step==8'h6f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1539[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1515[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1023[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1575[9:0] );

									end
									else
									if((r_sys_run_step==8'h65) || (r_sys_run_step==8'h67)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1443[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1311[9:0] );

									end
									else
									if((r_sys_run_step==8'h64) || (r_sys_run_step==8'h66)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1431[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1503[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp747[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp399[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp951[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1119[9:0] );

									end
									else
									if((r_sys_run_step==8'h45) || (r_sys_run_step==8'h47)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1059[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp687[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp291[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2079[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1875[9:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1779[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp471[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1707[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp267[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1047[9:0] );

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2055[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp387[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h3f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp963[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp759[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp303[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1203[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1299[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1671[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp279[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1491[9:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hb)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2241[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2553[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2133[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2121[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2565[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2145[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2361[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2289[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2181[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2541[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2469[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2253[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2169[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2193[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2157[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2349[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2445[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2337[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2457[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2529[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2265[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2325[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2229[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2421[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2517[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2109[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2385[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2373[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2277[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2481[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2433[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (8'h1c<=r_sys_run_step && r_sys_run_step<=8'h20)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (8'h1c<=r_sys_run_step && r_sys_run_step<=8'h20)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9b)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h26)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp41[9:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h93) || (r_sys_run_step==8'h95)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1995[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d) || (r_sys_run_step==8'h2f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp771[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp507[9:0] );

									end
									else
									if((r_sys_run_step==8'h94) || (r_sys_run_step==8'h96)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2007[9:0] );

									end
									else
									if((r_sys_run_step==8'h84) || (r_sys_run_step==8'h86)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1815[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1131[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp831[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp663[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1983[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1959[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp459[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp591[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp351[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1647[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1767[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp255[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1179[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1407[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1323[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1335[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1635[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1419[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1587[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1899[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e) || (r_sys_run_step==8'h30)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp783[9:0] );

									end
									else
									if((r_sys_run_step==8'h46) || (r_sys_run_step==8'h48)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1071[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1155[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1599[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e) || (r_sys_run_step==8'h40)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp975[9:0] );

									end
									else
									if((r_sys_run_step==8'h83) || (r_sys_run_step==8'h85)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1803[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp447[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1971[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp567[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1035[9:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1755[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1383[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1695[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp495[9:0] );

									end
									else
									if((r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1911[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp711[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp723[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp363[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp603[9:0] );

									end
									else
									if((r_sys_run_step==8'h55) || (r_sys_run_step==8'h57)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1251[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp543[9:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp855[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp699[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1287[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1107[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp819[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1167[9:0] );

									end
									else
									if((r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1719[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1851[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp651[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp483[9:0] );

									end
									else
									if((r_sys_run_step==8'h36) || (r_sys_run_step==8'h38)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp879[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp843[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp675[9:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1215[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp375[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp579[9:0] );

									end
									else
									if((r_sys_run_step==8'h54) || (r_sys_run_step==8'h56)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1239[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1863[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2067[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1611[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp555[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1011[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1659[9:0] );

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2043[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1395[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp639[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1227[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1623[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp735[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1191[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp315[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2091[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp915[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1479[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp231[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1527[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1683[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1143[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp411[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1791[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp243[9:0] );

									end
									else
									if((r_sys_run_step==8'h35) || (r_sys_run_step==8'h37)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp867[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1947[9:0] );

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1887[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d) || (r_sys_run_step==8'h5f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1347[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp939[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp927[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d) || (r_sys_run_step==8'h6f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1539[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1515[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1023[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1575[9:0] );

									end
									else
									if((r_sys_run_step==8'h65) || (r_sys_run_step==8'h67)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1443[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1311[9:0] );

									end
									else
									if((r_sys_run_step==8'h64) || (r_sys_run_step==8'h66)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1431[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1503[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp747[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp399[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp951[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1119[9:0] );

									end
									else
									if((r_sys_run_step==8'h45) || (r_sys_run_step==8'h47)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1059[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp687[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp291[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2079[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1875[9:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1779[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp471[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1707[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp267[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1047[9:0] );

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2055[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp387[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h3f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp963[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp759[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp303[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1203[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1299[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1671[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp279[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1491[9:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hb)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2241[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2553[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2133[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2121[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2565[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2145[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2361[9:0] );

									end
									else
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h11)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2289[9:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2181[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2541[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2469[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2253[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2169[9:0] );

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2193[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2157[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2349[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2445[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2337[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2457[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2529[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2265[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2325[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2229[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2421[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2517[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2109[9:0] );

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2385[9:0] );

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h18)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2373[9:0] );

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h10)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2277[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2481[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2433[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_V_3_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9b)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h26)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_V_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_tmp14;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_run_k_29 <= w_sys_tmp2102;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_tmp2103;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_run_k_29 <= w_sys_tmp2576;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_run_k_29 <= w_sys_tmp2596;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h9d)) begin
										r_run_k_29 <= w_sys_tmp3673;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_tmp3674;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h28)) begin
										r_run_k_29 <= w_sys_tmp3913;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_tmp3914;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h75)) begin
										r_run_k_29 <= w_sys_tmp4505;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_29 <= w_sys_tmp4506;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_run_k_29 <= w_sys_tmp4662;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_30 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_run_j_30 <= w_sys_tmp48;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_30 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h2) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc)) begin
										r_run_j_30 <= w_sys_tmp2611;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_run_j_30 <= w_sys_tmp2684;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_run_j_30 <= w_sys_tmp2696;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_n_31 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_n_31 <= w_sys_tmp2579;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_mx_32 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_my_33 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dt_34 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dx_35 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dy_36 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r1_37 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r2_38 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r3_39 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r4_40 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h10) || (r_sys_run_step==8'h11)) begin
										r_run_YY_41 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14)) begin
										r_run_YY_41 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_kx_42 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_ky_43 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_nlast_44 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_45 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_run_copy0_j_45 <= w_sys_tmp45;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy1_j_46 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (8'h1c<=r_sys_run_step && r_sys_run_step<=8'h20)) begin
										r_run_copy1_j_46 <= w_sys_tmp46;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy2_j_47 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_run_copy2_j_47 <= w_sys_tmp47;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_48 <= r_run_j_30;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd)) begin
										r_run_copy0_j_48 <= w_sys_tmp2610;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h98)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3626[9:0] );

									end
									else
									if((r_sys_run_step==8'h9c)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3662[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3656[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3650[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3644[9:0] );

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3620[9:0] );

									end
									else
									if((r_sys_run_step==8'h9d)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp3668[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h97)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp1995[9:0] );

									end
									else
									if((r_sys_run_step==8'h9c)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2079[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2067[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2055[9:0] );

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2007[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2043[9:0] );

									end
									else
									if((r_sys_run_step==8'h9d)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp2091[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h97)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp1995[9:0] );

									end
									else
									if((r_sys_run_step==8'h9c)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2079[9:0] );

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2067[9:0] );

									end
									else
									if((r_sys_run_step==8'h9a)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2055[9:0] );

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2007[9:0] );

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2043[9:0] );

									end
									else
									if((r_sys_run_step==8'h9d)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp2091[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h97<=r_sys_run_step && r_sys_run_step<=8'h9d)) begin
										r_sub19_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4486[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4491[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4501[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4496[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4481[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4f)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3200[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3194[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3152[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3176[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3188[9:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3182[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp3158[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4c)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1119[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1107[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1059[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1143[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1131[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1155[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp1071[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4c)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1119[9:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1107[9:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1059[9:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1143[9:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1131[9:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1155[9:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp1071[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h49<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sub09_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4196[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4201[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4191[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4211[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4206[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h43)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3128[9:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3140[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3104[9:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3152[9:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3134[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3110[9:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3146[9:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp3158[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h44)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1023[9:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1059[9:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1035[9:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1047[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp963[9:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1071[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp975[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1011[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h44)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1023[9:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1059[9:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1035[9:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1047[9:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp963[9:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1071[9:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp975[9:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1011[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h41<=r_sys_run_step && r_sys_run_step<=8'h48)) begin
										r_sub08_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4176[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4186[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4181[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4161[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4166[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp4171[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub24_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub24_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3890[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3860[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3902[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3908[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3884[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3896[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp3866[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_T_datain <= w_sys_tmp3682;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h26)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2541[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2469[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2553[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2529[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2565[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2481[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp2517[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_V_datain <= w_sys_tmp2117;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h26)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2541[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2469[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2553[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2529[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2565[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2481[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp2517[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_U_datain <= w_sys_tmp2111;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub24_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp4658[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp4653[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp4643[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp4638[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp4648[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub22_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub22_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3812[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3764[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3806[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3818[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3794[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3800[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3788[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp3770[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_T_datain <= w_sys_tmp3682;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2349[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2337[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2385[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2373[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2325[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2277[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2361[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp2289[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_V_datain <= w_sys_tmp2117;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2349[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2337[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2385[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2373[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2325[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2277[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2361[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp2289[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_U_datain <= w_sys_tmp2111;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub22_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4603[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4588[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4598[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4583[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4578[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp4593[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub23_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub23_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3812[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3860[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3848[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3818[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3842[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3836[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3866[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp3854[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_T_datain <= w_sys_tmp3682;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2445[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2469[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2457[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2385[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2373[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2421[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2481[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp2433[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_V_datain <= w_sys_tmp2117;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2445[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2469[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2457[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2385[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2373[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2421[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2481[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp2433[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_U_datain <= w_sys_tmp2111;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub23_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4618[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4633[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4608[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4628[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4613[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp4623[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h60)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3290[9:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3332[9:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3326[9:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3338[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3296[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3320[9:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3344[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp3314[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h65)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1419[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1383[9:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1431[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1347[9:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1443[9:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1407[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1395[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp1335[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h65)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1419[9:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1383[9:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1431[9:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1347[9:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1443[9:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1407[9:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1395[9:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp1335[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h60<=r_sys_run_step && r_sys_run_step<=8'h67)) begin
										r_sub12_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4286[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4296[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4291[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4281[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4301[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp4276[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2870[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2876[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2900[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2918[9:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2912[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2906[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2924[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp2894[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1f)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp579[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp567[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp591[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp603[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp507[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp495[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp543[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp555[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1f)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp579[9:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp567[9:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp591[9:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp603[9:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp507[9:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp495[9:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp543[9:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp555[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h1a<=r_sys_run_step && r_sys_run_step<=8'h21)) begin
										r_sub03_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4031[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4041[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4036[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4026[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4021[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4016[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2870[9:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2852[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2822[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2876[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2846[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2828[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2864[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp2858[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp459[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp507[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp495[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp411[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp471[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp483[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp447[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp399[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp459[9:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp507[9:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp495[9:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp411[9:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp471[9:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp483[9:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp447[9:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp399[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h12<=r_sys_run_step && r_sys_run_step<=8'h19)) begin
										r_sub02_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3991[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp4011[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3986[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp4006[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp4001[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3996[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5e)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3290[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3272[9:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3242[9:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3296[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3266[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3284[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3278[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp3248[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h58)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1239[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1311[9:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1347[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1251[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1299[9:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1335[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1323[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp1287[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h58)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1239[9:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1311[9:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1347[9:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1251[9:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1299[9:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1335[9:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1323[9:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp1287[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h58<=r_sys_run_step && r_sys_run_step<=8'h5f)) begin
										r_sub11_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4271[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4261[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4256[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4266[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4251[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4246[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h75)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3428[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3434[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3422[9:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3416[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3392[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3410[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3386[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h73)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1587[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1575[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1527[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1611[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1623[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1539[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp1599[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h73)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1587[9:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1575[9:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1527[9:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1611[9:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1623[9:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1539[9:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp1599[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h70<=r_sys_run_step && r_sys_run_step<=8'h76)) begin
										r_sub14_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4356[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4351[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4336[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4341[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4346[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h10)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2822[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2804[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2828[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2774[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2798[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2816[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2780[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp2810[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'he)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp375[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp363[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp351[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp387[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp411[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp303[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp315[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp399[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'he)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp375[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp363[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp351[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp387[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp411[9:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp303[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp315[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp399[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub01_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3956[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3971[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3966[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3961[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3981[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3976[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2738[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2768[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2762[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2774[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2780[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2750[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2744[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp2756[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp231[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp267[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp291[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp255[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp303[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp315[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp279[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp243[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp231[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp267[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp291[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp255[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp303[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp315[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp279[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp243[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub00_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3926[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3932[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3938[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3944[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3950[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3920[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6b)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3368[9:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3392[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3338[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3380[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3374[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3362[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3344[9:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3386[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6e)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1527[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1431[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1503[9:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1539[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1443[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1515[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1491[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp1479[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6e)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1527[9:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1431[9:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1503[9:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1539[9:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1443[9:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1515[9:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1491[9:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp1479[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h68<=r_sys_run_step && r_sys_run_step<=8'h6f)) begin
										r_sub13_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4331[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4326[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4321[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4311[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4316[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4306[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3d)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3092[9:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3104[9:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3110[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3098[9:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3056[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3086[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3062[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp3080[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h39)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp867[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp939[9:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp963[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp927[9:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp975[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp915[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp879[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp951[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h39)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp867[9:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp939[9:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp963[9:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp927[9:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp975[9:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp915[9:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp879[9:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp951[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h39<=r_sys_run_step && r_sys_run_step<=8'h40)) begin
										r_sub07_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4156[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4131[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4151[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4146[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4141[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp4136[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h85)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3524[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3506[9:0] );

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3512[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3482[9:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3476[9:0] );

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3530[9:0] );

									end
									else
									if((r_sys_run_step==8'h84)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3518[9:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3500[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7f)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1707[9:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1755[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1719[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1767[9:0] );

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1815[9:0] );

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1779[9:0] );

									end
									else
									if((r_sys_run_step==8'h84)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1791[9:0] );

									end
									else
									if((r_sys_run_step==8'h85)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp1803[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7f)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1707[9:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1755[9:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1719[9:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1767[9:0] );

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1815[9:0] );

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1779[9:0] );

									end
									else
									if((r_sys_run_step==8'h84)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1791[9:0] );

									end
									else
									if((r_sys_run_step==8'h85)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp1803[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h7f<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_sub16_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4406[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4401[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4411[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4396[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4391[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp4416[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h35)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3044[9:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3038[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3008[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3014[9:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3056[9:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3062[9:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3050[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp3032[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h37)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp867[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp771[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp819[9:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp831[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp783[9:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp855[9:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp879[9:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp843[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h37)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp867[9:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp771[9:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp819[9:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp831[9:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp783[9:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp855[9:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp879[9:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp843[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h31<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_sub06_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4101[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4126[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4121[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4106[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4116[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4111[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h78)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3446[9:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3482[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3464[9:0] );

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3476[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3440[9:0] );

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3470[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3452[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3458[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7d)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1707[9:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1719[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1659[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1683[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1647[9:0] );

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1695[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1671[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp1635[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7d)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1707[9:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1719[9:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1659[9:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1683[9:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1647[9:0] );

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1695[9:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1671[9:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp1635[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h77<=r_sys_run_step && r_sys_run_step<=8'h7e)) begin
										r_sub15_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4386[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4361[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4381[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4376[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4371[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp4366[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2e)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp3002[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2978[9:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2984[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2990[9:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp3008[9:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp3014[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2996[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2972[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2b)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp723[9:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp771[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp759[9:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp783[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp747[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp735[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp711[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp699[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2b)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp723[9:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp771[9:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp759[9:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp783[9:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp747[9:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp735[9:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp711[9:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp699[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h29<=r_sys_run_step && r_sys_run_step<=8'h30)) begin
										r_sub05_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4081[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4086[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4071[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4096[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4091[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4076[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h93)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3608[9:0] );

									end
									else
									if((r_sys_run_step==8'h96)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3626[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3578[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3602[9:0] );

									end
									else
									if((r_sys_run_step==8'h94)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3614[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3596[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3572[9:0] );

									end
									else
									if((r_sys_run_step==8'h95)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp3620[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h94)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1983[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1959[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1947[9:0] );

									end
									else
									if((r_sys_run_step==8'h95)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1995[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1899[9:0] );

									end
									else
									if((r_sys_run_step==8'h96)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp2007[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1911[9:0] );

									end
									else
									if((r_sys_run_step==8'h93)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp1971[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h94)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1983[9:0] );

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1959[9:0] );

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1947[9:0] );

									end
									else
									if((r_sys_run_step==8'h95)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1995[9:0] );

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1899[9:0] );

									end
									else
									if((r_sys_run_step==8'h96)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp2007[9:0] );

									end
									else
									if((r_sys_run_step==8'h90)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1911[9:0] );

									end
									else
									if((r_sys_run_step==8'h93)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp1971[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h8f<=r_sys_run_step && r_sys_run_step<=8'h96)) begin
										r_sub18_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4451[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4456[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4471[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4476[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4461[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4466[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h27)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2960[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2948[9:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2942[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2966[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2918[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2924[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp2954[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h24)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp639[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp591[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp687[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp603[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp651[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp675[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp663[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h24)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp639[9:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp591[9:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp687[9:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp603[9:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp651[9:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp675[9:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp663[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h22<=r_sys_run_step && r_sys_run_step<=8'h28)) begin
										r_sub04_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4066[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4051[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4056[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4061[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp4046[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h87)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3524[9:0] );

									end
									else
									if((r_sys_run_step==8'h8e)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3578[9:0] );

									end
									else
									if((r_sys_run_step==8'h8d)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3572[9:0] );

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3554[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3548[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3560[9:0] );

									end
									else
									if((r_sys_run_step==8'h8c)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3566[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3530[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8d)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1899[9:0] );

									end
									else
									if((r_sys_run_step==8'h8c)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1887[9:0] );

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1863[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1875[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1851[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1815[9:0] );

									end
									else
									if((r_sys_run_step==8'h8e)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1911[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp1803[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8d)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1899[9:0] );

									end
									else
									if((r_sys_run_step==8'h8c)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1887[9:0] );

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1863[9:0] );

									end
									else
									if((r_sys_run_step==8'h8b)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1875[9:0] );

									end
									else
									if((r_sys_run_step==8'h89)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1851[9:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1815[9:0] );

									end
									else
									if((r_sys_run_step==8'h8e)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1911[9:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp1803[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h87<=r_sys_run_step && r_sys_run_step<=8'h8e)) begin
										r_sub17_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4431[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4436[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4421[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4441[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4446[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp4426[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h52)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3218[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3212[9:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3242[9:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3236[9:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3230[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3206[9:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3248[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp3224[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_T_datain <= w_sys_tmp2740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h56)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1239[9:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1227[9:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1251[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1167[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1203[9:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1191[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1179[9:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp1215[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_V_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h56)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1239[9:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1227[9:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1251[9:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1167[9:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1203[9:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1191[9:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1179[9:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp1215[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_U_datain <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h50<=r_sys_run_step && r_sys_run_step<=8'h57)) begin
										r_sub10_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4236[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4226[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4241[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4221[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4231[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4216[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub20_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub20_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3698[9:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3716[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3722[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3680[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3686[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3710[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3692[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp3704[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_T_datain <= w_sys_tmp3682;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2181[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2157[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2169[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2133[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2121[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2145[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2193[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp2109[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_V_datain <= w_sys_tmp2117;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2181[9:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2157[9:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2169[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2133[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2121[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2145[9:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2193[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp2109[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_U_datain <= w_sys_tmp2111;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h9)) begin
										r_sub20_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4542[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4536[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4524[9:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4512[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4530[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp4518[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub21_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub21_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3716[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3764[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3722[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3758[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3740[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3746[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3752[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp3770[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_T_datain <= w_sys_tmp3682;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2181[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2253[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2241[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2265[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2277[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2229[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2193[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp2289[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_V_datain <= w_sys_tmp2117;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2181[9:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2253[9:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2241[9:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2265[9:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2277[9:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2229[9:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2193[9:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp2289[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_U_datain <= w_sys_tmp2111;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'ha<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_sub21_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4548[9:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4568[9:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4553[9:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4563[9:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4558[9:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp4573[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp0_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp1_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h19)) begin
										r_sys_tmp2_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp2_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h17)) begin
										r_sys_tmp3_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp3_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'hd)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp4_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp5_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp5_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp6_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp6_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp7_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp7_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp8_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp8_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp9_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp9_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp10_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp10_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp11_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp11_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp12_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp12_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp13_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp13_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp14_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp14_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp15_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp15_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp16_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp16_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp17_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp17_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp18_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp18_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp19_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp19_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp20_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp20_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp21_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp21_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp22_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp22_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp23_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp23_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp24_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp24_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp25_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp25_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp26_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp26_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp27_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp27_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp28_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp29_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp30_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp31_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp32_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp33_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp34_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp35_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp36_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp37_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp38_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp39_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp40_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp41_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp42_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp43_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp44_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp45_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp46_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp47_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp48_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp49_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp50_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp51_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp52_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp53_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp54_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp55_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp56_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp57_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp58_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp59_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp60_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp61_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp62_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp63_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp64_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp65_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp66_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp67_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp68_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp69_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp70_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp71_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp72_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp73_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp74_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp75_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp76_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp77_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp78_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp79_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp80_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp81_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp82_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp83_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp84_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp85_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp86_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp87_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp88_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp89_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp90_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp91_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp92_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp93_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp94_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp95_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp96_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp97_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp98_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp99_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp100_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp101_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp102_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp103_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp104_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp105_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp106_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp107_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp108_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp109_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
