/*
TimeStamp:	2016/5/10		14:45
*/


module c1_test03(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 5:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 5:0] w_sys_run_step_p1;
	wire signed [ 9:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [ 9:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [ 9:0] w_fld_uu_1_addr_0;
	wire        [31:0] w_fld_uu_1_datain_0;
	wire        [31:0] w_fld_uu_1_dataout_0;
	wire               w_fld_uu_1_r_w_0;
	wire               w_fld_uu_1_ce_0;
	reg  signed [ 9:0] r_fld_uu_1_addr_1;
	reg         [31:0] r_fld_uu_1_datain_1;
	wire        [31:0] w_fld_uu_1_dataout_1;
	reg                r_fld_uu_1_r_w_1;
	wire               w_fld_uu_1_ce_1;
	reg  signed [31:0] r_run_k_18;
	reg  signed [31:0] r_run_j_19;
	reg  signed [31:0] r_run_n_20;
	reg  signed [31:0] r_run_mx_21;
	reg  signed [31:0] r_run_my_22;
	reg  signed [31:0] r_run_nlast_23;
	reg  signed [31:0] r_run_copy0_j_24;
	reg  signed [31:0] r_run_copy0_j_25;
	reg  signed [31:0] r_run_copy1_j_26;
	reg  signed [31:0] r_run_copy2_j_27;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [ 9:0] w_sub09_u_addr;
	reg  signed [ 9:0] r_sub09_u_addr;
	wire        [31:0] w_sub09_u_datain;
	reg         [31:0] r_sub09_u_datain;
	wire        [31:0] w_sub09_u_dataout;
	wire               w_sub09_u_r_w;
	reg                r_sub09_u_r_w;
	wire signed [ 9:0] w_sub09_result_addr;
	reg  signed [ 9:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [ 9:0] w_sub08_u_addr;
	reg  signed [ 9:0] r_sub08_u_addr;
	wire        [31:0] w_sub08_u_datain;
	reg         [31:0] r_sub08_u_datain;
	wire        [31:0] w_sub08_u_dataout;
	wire               w_sub08_u_r_w;
	reg                r_sub08_u_r_w;
	wire signed [ 9:0] w_sub08_result_addr;
	reg  signed [ 9:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [ 9:0] w_sub12_u_addr;
	reg  signed [ 9:0] r_sub12_u_addr;
	wire        [31:0] w_sub12_u_datain;
	reg         [31:0] r_sub12_u_datain;
	wire        [31:0] w_sub12_u_dataout;
	wire               w_sub12_u_r_w;
	reg                r_sub12_u_r_w;
	wire signed [ 9:0] w_sub12_result_addr;
	reg  signed [ 9:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 9:0] w_sub03_u_addr;
	reg  signed [ 9:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [ 9:0] w_sub03_result_addr;
	reg  signed [ 9:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 9:0] w_sub02_u_addr;
	reg  signed [ 9:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [ 9:0] w_sub02_result_addr;
	reg  signed [ 9:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [ 9:0] w_sub11_u_addr;
	reg  signed [ 9:0] r_sub11_u_addr;
	wire        [31:0] w_sub11_u_datain;
	reg         [31:0] r_sub11_u_datain;
	wire        [31:0] w_sub11_u_dataout;
	wire               w_sub11_u_r_w;
	reg                r_sub11_u_r_w;
	wire signed [ 9:0] w_sub11_result_addr;
	reg  signed [ 9:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [ 9:0] w_sub14_u_addr;
	reg  signed [ 9:0] r_sub14_u_addr;
	wire        [31:0] w_sub14_u_datain;
	reg         [31:0] r_sub14_u_datain;
	wire        [31:0] w_sub14_u_dataout;
	wire               w_sub14_u_r_w;
	reg                r_sub14_u_r_w;
	wire signed [ 9:0] w_sub14_result_addr;
	reg  signed [ 9:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 9:0] w_sub01_u_addr;
	reg  signed [ 9:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [ 9:0] w_sub01_result_addr;
	reg  signed [ 9:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [ 9:0] w_sub13_u_addr;
	reg  signed [ 9:0] r_sub13_u_addr;
	wire        [31:0] w_sub13_u_datain;
	reg         [31:0] r_sub13_u_datain;
	wire        [31:0] w_sub13_u_dataout;
	wire               w_sub13_u_r_w;
	reg                r_sub13_u_r_w;
	wire signed [ 9:0] w_sub13_result_addr;
	reg  signed [ 9:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 9:0] w_sub00_u_addr;
	reg  signed [ 9:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [ 9:0] w_sub00_result_addr;
	reg  signed [ 9:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [ 9:0] w_sub07_u_addr;
	reg  signed [ 9:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [ 9:0] w_sub07_result_addr;
	reg  signed [ 9:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [ 9:0] w_sub06_u_addr;
	reg  signed [ 9:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [ 9:0] w_sub06_result_addr;
	reg  signed [ 9:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [ 9:0] w_sub15_u_addr;
	reg  signed [ 9:0] r_sub15_u_addr;
	wire        [31:0] w_sub15_u_datain;
	reg         [31:0] r_sub15_u_datain;
	wire        [31:0] w_sub15_u_dataout;
	wire               w_sub15_u_r_w;
	reg                r_sub15_u_r_w;
	wire signed [ 9:0] w_sub15_result_addr;
	reg  signed [ 9:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [ 9:0] w_sub05_u_addr;
	reg  signed [ 9:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [ 9:0] w_sub05_result_addr;
	reg  signed [ 9:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [ 9:0] w_sub04_u_addr;
	reg  signed [ 9:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [ 9:0] w_sub04_result_addr;
	reg  signed [ 9:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [ 9:0] w_sub10_u_addr;
	reg  signed [ 9:0] r_sub10_u_addr;
	wire        [31:0] w_sub10_u_datain;
	reg         [31:0] r_sub10_u_datain;
	wire        [31:0] w_sub10_u_dataout;
	wire               w_sub10_u_r_w;
	reg                r_sub10_u_r_w;
	wire signed [ 9:0] w_sub10_result_addr;
	reg  signed [ 9:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire               w_sys_tmp4;
	wire               w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire               w_sys_tmp7;
	wire               w_sys_tmp8;
	wire signed [31:0] w_sys_tmp11;
	wire signed [31:0] w_sys_tmp12;
	wire signed [31:0] w_sys_tmp13;
	wire        [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire               w_sys_tmp94;
	wire               w_sys_tmp95;
	wire signed [31:0] w_sys_tmp96;
	wire               w_sys_tmp97;
	wire               w_sys_tmp98;
	wire signed [31:0] w_sys_tmp101;
	wire signed [31:0] w_sys_tmp102;
	wire        [31:0] w_sys_tmp103;
	wire signed [31:0] w_sys_tmp105;
	wire signed [31:0] w_sys_tmp106;
	wire        [31:0] w_sys_tmp108;
	wire signed [31:0] w_sys_tmp110;
	wire signed [31:0] w_sys_tmp111;
	wire        [31:0] w_sys_tmp113;
	wire signed [31:0] w_sys_tmp115;
	wire signed [31:0] w_sys_tmp116;
	wire signed [31:0] w_sys_tmp119;
	wire signed [31:0] w_sys_tmp120;
	wire signed [31:0] w_sys_tmp121;
	wire signed [31:0] w_sys_tmp122;
	wire               w_sys_tmp261;
	wire               w_sys_tmp262;
	wire signed [31:0] w_sys_tmp263;
	wire signed [31:0] w_sys_tmp266;
	wire signed [31:0] w_sys_tmp267;
	wire        [31:0] w_sys_tmp268;
	wire signed [31:0] w_sys_tmp272;
	wire signed [31:0] w_sys_tmp273;
	wire signed [31:0] w_sys_tmp278;
	wire signed [31:0] w_sys_tmp279;
	wire signed [31:0] w_sys_tmp284;
	wire signed [31:0] w_sys_tmp285;
	wire signed [31:0] w_sys_tmp302;
	wire signed [31:0] w_sys_tmp303;
	wire signed [31:0] w_sys_tmp308;
	wire signed [31:0] w_sys_tmp309;
	wire signed [31:0] w_sys_tmp326;
	wire signed [31:0] w_sys_tmp327;
	wire signed [31:0] w_sys_tmp332;
	wire signed [31:0] w_sys_tmp333;
	wire signed [31:0] w_sys_tmp350;
	wire signed [31:0] w_sys_tmp351;
	wire signed [31:0] w_sys_tmp356;
	wire signed [31:0] w_sys_tmp357;
	wire signed [31:0] w_sys_tmp362;
	wire signed [31:0] w_sys_tmp363;
	wire signed [31:0] w_sys_tmp368;
	wire signed [31:0] w_sys_tmp369;
	wire signed [31:0] w_sys_tmp374;
	wire signed [31:0] w_sys_tmp375;
	wire signed [31:0] w_sys_tmp380;
	wire signed [31:0] w_sys_tmp381;
	wire signed [31:0] w_sys_tmp386;
	wire signed [31:0] w_sys_tmp387;
	wire signed [31:0] w_sys_tmp404;
	wire signed [31:0] w_sys_tmp405;
	wire signed [31:0] w_sys_tmp410;
	wire signed [31:0] w_sys_tmp411;
	wire signed [31:0] w_sys_tmp428;
	wire signed [31:0] w_sys_tmp429;
	wire signed [31:0] w_sys_tmp434;
	wire signed [31:0] w_sys_tmp435;
	wire signed [31:0] w_sys_tmp452;
	wire signed [31:0] w_sys_tmp453;
	wire signed [31:0] w_sys_tmp458;
	wire signed [31:0] w_sys_tmp459;
	wire signed [31:0] w_sys_tmp464;
	wire signed [31:0] w_sys_tmp465;
	wire signed [31:0] w_sys_tmp470;
	wire signed [31:0] w_sys_tmp471;
	wire signed [31:0] w_sys_tmp476;
	wire signed [31:0] w_sys_tmp477;
	wire signed [31:0] w_sys_tmp482;
	wire signed [31:0] w_sys_tmp483;
	wire signed [31:0] w_sys_tmp488;
	wire signed [31:0] w_sys_tmp489;
	wire signed [31:0] w_sys_tmp506;
	wire signed [31:0] w_sys_tmp507;
	wire signed [31:0] w_sys_tmp512;
	wire signed [31:0] w_sys_tmp513;
	wire signed [31:0] w_sys_tmp530;
	wire signed [31:0] w_sys_tmp531;
	wire signed [31:0] w_sys_tmp536;
	wire signed [31:0] w_sys_tmp537;
	wire signed [31:0] w_sys_tmp554;
	wire signed [31:0] w_sys_tmp555;
	wire signed [31:0] w_sys_tmp560;
	wire signed [31:0] w_sys_tmp561;
	wire signed [31:0] w_sys_tmp566;
	wire signed [31:0] w_sys_tmp567;
	wire signed [31:0] w_sys_tmp571;
	wire signed [31:0] w_sys_tmp572;
	wire               w_sys_tmp573;
	wire               w_sys_tmp574;
	wire signed [31:0] w_sys_tmp575;
	wire signed [31:0] w_sys_tmp578;
	wire signed [31:0] w_sys_tmp579;
	wire        [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp584;
	wire signed [31:0] w_sys_tmp585;
	wire signed [31:0] w_sys_tmp590;
	wire signed [31:0] w_sys_tmp591;
	wire signed [31:0] w_sys_tmp596;
	wire signed [31:0] w_sys_tmp597;
	wire signed [31:0] w_sys_tmp614;
	wire signed [31:0] w_sys_tmp615;
	wire signed [31:0] w_sys_tmp620;
	wire signed [31:0] w_sys_tmp621;
	wire signed [31:0] w_sys_tmp638;
	wire signed [31:0] w_sys_tmp639;
	wire signed [31:0] w_sys_tmp644;
	wire signed [31:0] w_sys_tmp645;
	wire signed [31:0] w_sys_tmp662;
	wire signed [31:0] w_sys_tmp663;
	wire signed [31:0] w_sys_tmp668;
	wire signed [31:0] w_sys_tmp669;
	wire signed [31:0] w_sys_tmp674;
	wire signed [31:0] w_sys_tmp675;
	wire signed [31:0] w_sys_tmp679;
	wire signed [31:0] w_sys_tmp680;
	wire               w_sys_tmp681;
	wire               w_sys_tmp682;
	wire signed [31:0] w_sys_tmp683;
	wire signed [31:0] w_sys_tmp686;
	wire signed [31:0] w_sys_tmp687;
	wire        [31:0] w_sys_tmp688;
	wire signed [31:0] w_sys_tmp692;
	wire signed [31:0] w_sys_tmp693;
	wire signed [31:0] w_sys_tmp698;
	wire signed [31:0] w_sys_tmp699;
	wire signed [31:0] w_sys_tmp703;
	wire signed [31:0] w_sys_tmp704;
	wire signed [31:0] w_sys_tmp708;
	wire signed [31:0] w_sys_tmp709;
	wire signed [31:0] w_sys_tmp713;
	wire signed [31:0] w_sys_tmp714;
	wire signed [31:0] w_sys_tmp718;
	wire signed [31:0] w_sys_tmp719;
	wire signed [31:0] w_sys_tmp723;
	wire signed [31:0] w_sys_tmp724;
	wire signed [31:0] w_sys_tmp728;
	wire signed [31:0] w_sys_tmp729;
	wire signed [31:0] w_sys_tmp733;
	wire signed [31:0] w_sys_tmp734;
	wire signed [31:0] w_sys_tmp738;
	wire signed [31:0] w_sys_tmp739;
	wire signed [31:0] w_sys_tmp743;
	wire signed [31:0] w_sys_tmp744;
	wire signed [31:0] w_sys_tmp748;
	wire signed [31:0] w_sys_tmp749;
	wire signed [31:0] w_sys_tmp753;
	wire signed [31:0] w_sys_tmp754;
	wire signed [31:0] w_sys_tmp758;
	wire signed [31:0] w_sys_tmp759;
	wire signed [31:0] w_sys_tmp763;
	wire signed [31:0] w_sys_tmp764;
	wire signed [31:0] w_sys_tmp768;
	wire signed [31:0] w_sys_tmp769;
	wire signed [31:0] w_sys_tmp773;
	wire signed [31:0] w_sys_tmp774;
	wire signed [31:0] w_sys_tmp778;
	wire signed [31:0] w_sys_tmp779;
	wire signed [31:0] w_sys_tmp783;
	wire signed [31:0] w_sys_tmp784;
	wire signed [31:0] w_sys_tmp788;
	wire signed [31:0] w_sys_tmp789;
	wire signed [31:0] w_sys_tmp793;
	wire signed [31:0] w_sys_tmp794;
	wire signed [31:0] w_sys_tmp798;
	wire signed [31:0] w_sys_tmp799;
	wire signed [31:0] w_sys_tmp803;
	wire signed [31:0] w_sys_tmp804;
	wire signed [31:0] w_sys_tmp808;
	wire signed [31:0] w_sys_tmp809;
	wire signed [31:0] w_sys_tmp813;
	wire signed [31:0] w_sys_tmp814;
	wire signed [31:0] w_sys_tmp818;
	wire signed [31:0] w_sys_tmp819;
	wire signed [31:0] w_sys_tmp822;
	wire signed [31:0] w_sys_tmp823;
	wire               w_sys_tmp824;
	wire               w_sys_tmp825;
	wire signed [31:0] w_sys_tmp826;
	wire signed [31:0] w_sys_tmp829;
	wire signed [31:0] w_sys_tmp830;
	wire        [31:0] w_sys_tmp831;
	wire signed [31:0] w_sys_tmp835;
	wire signed [31:0] w_sys_tmp836;
	wire signed [31:0] w_sys_tmp841;
	wire signed [31:0] w_sys_tmp842;
	wire signed [31:0] w_sys_tmp846;
	wire signed [31:0] w_sys_tmp847;
	wire signed [31:0] w_sys_tmp851;
	wire signed [31:0] w_sys_tmp852;
	wire signed [31:0] w_sys_tmp856;
	wire signed [31:0] w_sys_tmp857;
	wire signed [31:0] w_sys_tmp861;
	wire signed [31:0] w_sys_tmp862;
	wire signed [31:0] w_sys_tmp866;
	wire signed [31:0] w_sys_tmp867;
	wire signed [31:0] w_sys_tmp871;
	wire signed [31:0] w_sys_tmp872;
	wire signed [31:0] w_sys_tmp875;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 6'h1);
	assign w_fld_u_0_addr_0 = 10'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_fld_uu_1_addr_0 = 10'sh0;
	assign w_fld_uu_1_datain_0 = 32'h0;
	assign w_fld_uu_1_r_w_0 = 1'h0;
	assign w_fld_uu_1_ce_0 = w_sys_ce;
	assign w_fld_uu_1_ce_1 = w_sys_ce;
	assign w_sub09_u_addr = ( (|r_sys_processing_methodID) ? r_sub09_u_addr : 10'sh0 ) ;
	assign w_sub09_u_datain = ( (|r_sys_processing_methodID) ? r_sub09_u_datain : 32'h0 ) ;
	assign w_sub09_u_r_w = ( (|r_sys_processing_methodID) ? r_sub09_u_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 10'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_u_addr = ( (|r_sys_processing_methodID) ? r_sub08_u_addr : 10'sh0 ) ;
	assign w_sub08_u_datain = ( (|r_sys_processing_methodID) ? r_sub08_u_datain : 32'h0 ) ;
	assign w_sub08_u_r_w = ( (|r_sys_processing_methodID) ? r_sub08_u_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 10'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub12_u_addr = ( (|r_sys_processing_methodID) ? r_sub12_u_addr : 10'sh0 ) ;
	assign w_sub12_u_datain = ( (|r_sys_processing_methodID) ? r_sub12_u_datain : 32'h0 ) ;
	assign w_sub12_u_r_w = ( (|r_sys_processing_methodID) ? r_sub12_u_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 10'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 10'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 10'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 10'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 10'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_u_addr = ( (|r_sys_processing_methodID) ? r_sub11_u_addr : 10'sh0 ) ;
	assign w_sub11_u_datain = ( (|r_sys_processing_methodID) ? r_sub11_u_datain : 32'h0 ) ;
	assign w_sub11_u_r_w = ( (|r_sys_processing_methodID) ? r_sub11_u_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 10'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_u_addr = ( (|r_sys_processing_methodID) ? r_sub14_u_addr : 10'sh0 ) ;
	assign w_sub14_u_datain = ( (|r_sys_processing_methodID) ? r_sub14_u_datain : 32'h0 ) ;
	assign w_sub14_u_r_w = ( (|r_sys_processing_methodID) ? r_sub14_u_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 10'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 10'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 10'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub13_u_addr = ( (|r_sys_processing_methodID) ? r_sub13_u_addr : 10'sh0 ) ;
	assign w_sub13_u_datain = ( (|r_sys_processing_methodID) ? r_sub13_u_datain : 32'h0 ) ;
	assign w_sub13_u_r_w = ( (|r_sys_processing_methodID) ? r_sub13_u_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 10'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 10'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 10'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 10'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 10'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 10'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 10'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_u_addr = ( (|r_sys_processing_methodID) ? r_sub15_u_addr : 10'sh0 ) ;
	assign w_sub15_u_datain = ( (|r_sys_processing_methodID) ? r_sub15_u_datain : 32'h0 ) ;
	assign w_sub15_u_r_w = ( (|r_sys_processing_methodID) ? r_sub15_u_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 10'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 10'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 10'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 10'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 10'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_u_addr = ( (|r_sys_processing_methodID) ? r_sub10_u_addr : 10'sh0 ) ;
	assign w_sub10_u_datain = ( (|r_sys_processing_methodID) ? r_sub10_u_datain : 32'h0 ) ;
	assign w_sub10_u_r_w = ( (|r_sys_processing_methodID) ? r_sub10_u_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 10'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh0000000b;
	assign w_sys_tmp3 = 32'sh00000190;
	assign w_sys_tmp4 = ( !w_sys_tmp5 );
	assign w_sys_tmp5 = (r_run_my_22 < r_run_k_18);
	assign w_sys_tmp6 = (r_run_k_18 + w_sys_intOne);
	assign w_sys_tmp7 = ( !w_sys_tmp8 );
	assign w_sys_tmp8 = (r_run_mx_21 < r_run_j_19);
	assign w_sys_tmp11 = (w_sys_tmp12 + r_run_k_18);
	assign w_sys_tmp12 = (r_run_j_19 * w_sys_tmp13);
	assign w_sys_tmp13 = 32'sh0000000b;
	assign w_sys_tmp14 = 32'h0;
	assign w_sys_tmp16 = (w_sys_tmp17 + r_run_k_18);
	assign w_sys_tmp17 = (r_run_copy0_j_24 * w_sys_tmp13);
	assign w_sys_tmp20 = (r_run_copy0_j_24 + w_sys_intOne);
	assign w_sys_tmp21 = (r_run_j_19 + w_sys_intOne);
	assign w_sys_tmp94 = ( !w_sys_tmp95 );
	assign w_sys_tmp95 = (r_run_nlast_23 < r_run_n_20);
	assign w_sys_tmp96 = (r_run_n_20 + w_sys_intOne);
	assign w_sys_tmp97 = ( !w_sys_tmp98 );
	assign w_sys_tmp98 = (r_run_my_22 < r_run_j_19);
	assign w_sys_tmp101 = (w_sys_tmp102 + r_run_j_19);
	assign w_sys_tmp102 = 32'sh0000000b;
	assign w_sys_tmp103 = 32'h3f000000;
	assign w_sys_tmp105 = (w_sys_tmp106 + r_run_copy2_j_27);
	assign w_sys_tmp106 = (w_sys_tmp102 * r_run_mx_21);
	assign w_sys_tmp108 = 32'h0;
	assign w_sys_tmp110 = (w_sys_tmp111 + w_sys_intOne);
	assign w_sys_tmp111 = (r_run_copy1_j_26 * w_sys_tmp102);
	assign w_sys_tmp113 = 32'h3f800000;
	assign w_sys_tmp115 = (w_sys_tmp116 + r_run_my_22);
	assign w_sys_tmp116 = (r_run_copy0_j_25 * w_sys_tmp102);
	assign w_sys_tmp119 = (r_run_copy0_j_25 + w_sys_intOne);
	assign w_sys_tmp120 = (r_run_copy1_j_26 + w_sys_intOne);
	assign w_sys_tmp121 = (r_run_copy2_j_27 + w_sys_intOne);
	assign w_sys_tmp122 = (r_run_j_19 + w_sys_intOne);
	assign w_sys_tmp261 = ( !w_sys_tmp262 );
	assign w_sys_tmp262 = (w_sys_tmp263 < r_run_k_18);
	assign w_sys_tmp263 = 32'sh00000004;
	assign w_sys_tmp266 = (w_sys_tmp267 + r_run_k_18);
	assign w_sys_tmp267 = 32'sh0000000b;
	assign w_sys_tmp268 = w_fld_u_0_dataout_1;
	assign w_sys_tmp272 = (w_sys_tmp273 + r_run_k_18);
	assign w_sys_tmp273 = 32'sh00000016;
	assign w_sys_tmp278 = (w_sys_tmp279 + r_run_k_18);
	assign w_sys_tmp279 = 32'sh00000021;
	assign w_sys_tmp284 = (w_sys_tmp285 + r_run_k_18);
	assign w_sys_tmp285 = 32'sh0000002c;
	assign w_sys_tmp302 = (w_sys_tmp303 + r_run_k_18);
	assign w_sys_tmp303 = 32'sh00000037;
	assign w_sys_tmp308 = (w_sys_tmp309 + r_run_k_18);
	assign w_sys_tmp309 = 32'sh00000042;
	assign w_sys_tmp326 = (w_sys_tmp327 + r_run_k_18);
	assign w_sys_tmp327 = 32'sh0000004d;
	assign w_sys_tmp332 = (w_sys_tmp333 + r_run_k_18);
	assign w_sys_tmp333 = 32'sh00000058;
	assign w_sys_tmp350 = (w_sys_tmp351 + r_run_k_18);
	assign w_sys_tmp351 = 32'sh00000063;
	assign w_sys_tmp356 = (w_sys_tmp357 + r_run_k_18);
	assign w_sys_tmp357 = 32'sh0000006e;
	assign w_sys_tmp362 = (w_sys_tmp363 + r_run_k_18);
	assign w_sys_tmp363 = 32'sh00000079;
	assign w_sys_tmp368 = (w_sys_tmp369 + r_run_k_18);
	assign w_sys_tmp369 = 32'sh0000000d;
	assign w_sys_tmp374 = (w_sys_tmp375 + r_run_k_18);
	assign w_sys_tmp375 = 32'sh00000018;
	assign w_sys_tmp380 = (w_sys_tmp381 + r_run_k_18);
	assign w_sys_tmp381 = 32'sh00000023;
	assign w_sys_tmp386 = (w_sys_tmp387 + r_run_k_18);
	assign w_sys_tmp387 = 32'sh0000002e;
	assign w_sys_tmp404 = (w_sys_tmp405 + r_run_k_18);
	assign w_sys_tmp405 = 32'sh00000039;
	assign w_sys_tmp410 = (w_sys_tmp411 + r_run_k_18);
	assign w_sys_tmp411 = 32'sh00000044;
	assign w_sys_tmp428 = (w_sys_tmp429 + r_run_k_18);
	assign w_sys_tmp429 = 32'sh0000004f;
	assign w_sys_tmp434 = (w_sys_tmp435 + r_run_k_18);
	assign w_sys_tmp435 = 32'sh0000005a;
	assign w_sys_tmp452 = (w_sys_tmp453 + r_run_k_18);
	assign w_sys_tmp453 = 32'sh00000065;
	assign w_sys_tmp458 = (w_sys_tmp459 + r_run_k_18);
	assign w_sys_tmp459 = 32'sh00000070;
	assign w_sys_tmp464 = (w_sys_tmp465 + r_run_k_18);
	assign w_sys_tmp465 = 32'sh0000007b;
	assign w_sys_tmp470 = (w_sys_tmp471 + r_run_k_18);
	assign w_sys_tmp471 = 32'sh0000000f;
	assign w_sys_tmp476 = (w_sys_tmp477 + r_run_k_18);
	assign w_sys_tmp477 = 32'sh0000001a;
	assign w_sys_tmp482 = (w_sys_tmp483 + r_run_k_18);
	assign w_sys_tmp483 = 32'sh00000025;
	assign w_sys_tmp488 = (w_sys_tmp489 + r_run_k_18);
	assign w_sys_tmp489 = 32'sh00000030;
	assign w_sys_tmp506 = (w_sys_tmp507 + r_run_k_18);
	assign w_sys_tmp507 = 32'sh0000003b;
	assign w_sys_tmp512 = (w_sys_tmp513 + r_run_k_18);
	assign w_sys_tmp513 = 32'sh00000046;
	assign w_sys_tmp530 = (w_sys_tmp531 + r_run_k_18);
	assign w_sys_tmp531 = 32'sh00000051;
	assign w_sys_tmp536 = (w_sys_tmp537 + r_run_k_18);
	assign w_sys_tmp537 = 32'sh0000005c;
	assign w_sys_tmp554 = (w_sys_tmp555 + r_run_k_18);
	assign w_sys_tmp555 = 32'sh00000067;
	assign w_sys_tmp560 = (w_sys_tmp561 + r_run_k_18);
	assign w_sys_tmp561 = 32'sh00000072;
	assign w_sys_tmp566 = (w_sys_tmp567 + r_run_k_18);
	assign w_sys_tmp567 = 32'sh0000007d;
	assign w_sys_tmp571 = (r_run_k_18 + w_sys_intOne);
	assign w_sys_tmp572 = 32'sh00000007;
	assign w_sys_tmp573 = ( !w_sys_tmp574 );
	assign w_sys_tmp574 = (w_sys_tmp575 < r_run_k_18);
	assign w_sys_tmp575 = 32'sh0000000b;
	assign w_sys_tmp578 = (w_sys_tmp579 + r_run_k_18);
	assign w_sys_tmp579 = 32'sh0000000b;
	assign w_sys_tmp580 = w_fld_u_0_dataout_1;
	assign w_sys_tmp584 = (w_sys_tmp585 + r_run_k_18);
	assign w_sys_tmp585 = 32'sh00000016;
	assign w_sys_tmp590 = (w_sys_tmp591 + r_run_k_18);
	assign w_sys_tmp591 = 32'sh00000021;
	assign w_sys_tmp596 = (w_sys_tmp597 + r_run_k_18);
	assign w_sys_tmp597 = 32'sh0000002c;
	assign w_sys_tmp614 = (w_sys_tmp615 + r_run_k_18);
	assign w_sys_tmp615 = 32'sh00000037;
	assign w_sys_tmp620 = (w_sys_tmp621 + r_run_k_18);
	assign w_sys_tmp621 = 32'sh00000042;
	assign w_sys_tmp638 = (w_sys_tmp639 + r_run_k_18);
	assign w_sys_tmp639 = 32'sh0000004d;
	assign w_sys_tmp644 = (w_sys_tmp645 + r_run_k_18);
	assign w_sys_tmp645 = 32'sh00000058;
	assign w_sys_tmp662 = (w_sys_tmp663 + r_run_k_18);
	assign w_sys_tmp663 = 32'sh00000063;
	assign w_sys_tmp668 = (w_sys_tmp669 + r_run_k_18);
	assign w_sys_tmp669 = 32'sh0000006e;
	assign w_sys_tmp674 = (w_sys_tmp675 + r_run_k_18);
	assign w_sys_tmp675 = 32'sh00000079;
	assign w_sys_tmp679 = (r_run_k_18 + w_sys_intOne);
	assign w_sys_tmp680 = 32'sh00000002;
	assign w_sys_tmp681 = ( !w_sys_tmp682 );
	assign w_sys_tmp682 = (w_sys_tmp683 < r_run_k_18);
	assign w_sys_tmp683 = 32'sh00000003;
	assign w_sys_tmp686 = (w_sys_tmp687 + r_run_k_18);
	assign w_sys_tmp687 = 32'sh00000016;
	assign w_sys_tmp688 = w_sub00_result_dataout;
	assign w_sys_tmp692 = (w_sys_tmp693 + r_run_k_18);
	assign w_sys_tmp693 = 32'sh00000021;
	assign w_sys_tmp698 = (w_sys_tmp699 + r_run_k_18);
	assign w_sys_tmp699 = 32'sh0000002c;
	assign w_sys_tmp703 = (w_sys_tmp704 + r_run_k_18);
	assign w_sys_tmp704 = 32'sh00000037;
	assign w_sys_tmp708 = (w_sys_tmp709 + r_run_k_18);
	assign w_sys_tmp709 = 32'sh00000042;
	assign w_sys_tmp713 = (w_sys_tmp714 + r_run_k_18);
	assign w_sys_tmp714 = 32'sh0000004d;
	assign w_sys_tmp718 = (w_sys_tmp719 + r_run_k_18);
	assign w_sys_tmp719 = 32'sh00000058;
	assign w_sys_tmp723 = (w_sys_tmp724 + r_run_k_18);
	assign w_sys_tmp724 = 32'sh00000063;
	assign w_sys_tmp728 = (w_sys_tmp729 + r_run_k_18);
	assign w_sys_tmp729 = 32'sh0000006e;
	assign w_sys_tmp733 = (w_sys_tmp734 + r_run_k_18);
	assign w_sys_tmp734 = 32'sh00000018;
	assign w_sys_tmp738 = (w_sys_tmp739 + r_run_k_18);
	assign w_sys_tmp739 = 32'sh00000023;
	assign w_sys_tmp743 = (w_sys_tmp744 + r_run_k_18);
	assign w_sys_tmp744 = 32'sh0000002e;
	assign w_sys_tmp748 = (w_sys_tmp749 + r_run_k_18);
	assign w_sys_tmp749 = 32'sh00000039;
	assign w_sys_tmp753 = (w_sys_tmp754 + r_run_k_18);
	assign w_sys_tmp754 = 32'sh00000044;
	assign w_sys_tmp758 = (w_sys_tmp759 + r_run_k_18);
	assign w_sys_tmp759 = 32'sh0000004f;
	assign w_sys_tmp763 = (w_sys_tmp764 + r_run_k_18);
	assign w_sys_tmp764 = 32'sh0000005a;
	assign w_sys_tmp768 = (w_sys_tmp769 + r_run_k_18);
	assign w_sys_tmp769 = 32'sh00000065;
	assign w_sys_tmp773 = (w_sys_tmp774 + r_run_k_18);
	assign w_sys_tmp774 = 32'sh00000070;
	assign w_sys_tmp778 = (w_sys_tmp779 + r_run_k_18);
	assign w_sys_tmp779 = 32'sh0000001a;
	assign w_sys_tmp783 = (w_sys_tmp784 + r_run_k_18);
	assign w_sys_tmp784 = 32'sh00000025;
	assign w_sys_tmp788 = (w_sys_tmp789 + r_run_k_18);
	assign w_sys_tmp789 = 32'sh00000030;
	assign w_sys_tmp793 = (w_sys_tmp794 + r_run_k_18);
	assign w_sys_tmp794 = 32'sh0000003b;
	assign w_sys_tmp798 = (w_sys_tmp799 + r_run_k_18);
	assign w_sys_tmp799 = 32'sh00000046;
	assign w_sys_tmp803 = (w_sys_tmp804 + r_run_k_18);
	assign w_sys_tmp804 = 32'sh00000051;
	assign w_sys_tmp808 = (w_sys_tmp809 + r_run_k_18);
	assign w_sys_tmp809 = 32'sh0000005c;
	assign w_sys_tmp813 = (w_sys_tmp814 + r_run_k_18);
	assign w_sys_tmp814 = 32'sh00000067;
	assign w_sys_tmp818 = (w_sys_tmp819 + r_run_k_18);
	assign w_sys_tmp819 = 32'sh00000072;
	assign w_sys_tmp822 = (r_run_k_18 + w_sys_intOne);
	assign w_sys_tmp823 = 32'sh00000008;
	assign w_sys_tmp824 = ( !w_sys_tmp825 );
	assign w_sys_tmp825 = (w_sys_tmp826 < r_run_k_18);
	assign w_sys_tmp826 = 32'sh0000000a;
	assign w_sys_tmp829 = (w_sys_tmp830 + r_run_k_18);
	assign w_sys_tmp830 = 32'sh00000016;
	assign w_sys_tmp831 = w_sub12_result_dataout;
	assign w_sys_tmp835 = (w_sys_tmp836 + r_run_k_18);
	assign w_sys_tmp836 = 32'sh00000021;
	assign w_sys_tmp841 = (w_sys_tmp842 + r_run_k_18);
	assign w_sys_tmp842 = 32'sh0000002c;
	assign w_sys_tmp846 = (w_sys_tmp847 + r_run_k_18);
	assign w_sys_tmp847 = 32'sh00000037;
	assign w_sys_tmp851 = (w_sys_tmp852 + r_run_k_18);
	assign w_sys_tmp852 = 32'sh00000042;
	assign w_sys_tmp856 = (w_sys_tmp857 + r_run_k_18);
	assign w_sys_tmp857 = 32'sh0000004d;
	assign w_sys_tmp861 = (w_sys_tmp862 + r_run_k_18);
	assign w_sys_tmp862 = 32'sh00000058;
	assign w_sys_tmp866 = (w_sys_tmp867 + r_run_k_18);
	assign w_sys_tmp867 = 32'sh00000063;
	assign w_sys_tmp871 = (w_sys_tmp872 + r_run_k_18);
	assign w_sys_tmp872 = 32'sh0000006e;
	assign w_sys_tmp875 = (r_run_k_18 + w_sys_intOne);


	sub09
		sub09_inst(
			.i_fld_result_1_addr_0 (w_sub09_result_addr),
			.i_fld_result_1_datain_0 (w_sub09_result_datain),
			.o_fld_result_1_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub09_result_r_w),
			.i_fld_u_0_addr_0 (w_sub09_u_addr),
			.i_fld_u_0_datain_0 (w_sub09_u_datain),
			.o_fld_u_0_dataout_0 (w_sub09_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub09_u_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_result_1_addr_0 (w_sub08_result_addr),
			.i_fld_result_1_datain_0 (w_sub08_result_datain),
			.o_fld_result_1_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub08_result_r_w),
			.i_fld_u_0_addr_0 (w_sub08_u_addr),
			.i_fld_u_0_datain_0 (w_sub08_u_datain),
			.o_fld_u_0_dataout_0 (w_sub08_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub08_u_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_result_1_addr_0 (w_sub12_result_addr),
			.i_fld_result_1_datain_0 (w_sub12_result_datain),
			.o_fld_result_1_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub12_result_r_w),
			.i_fld_u_0_addr_0 (w_sub12_u_addr),
			.i_fld_u_0_datain_0 (w_sub12_u_datain),
			.o_fld_u_0_dataout_0 (w_sub12_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub12_u_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_result_1_addr_0 (w_sub11_result_addr),
			.i_fld_result_1_datain_0 (w_sub11_result_datain),
			.o_fld_result_1_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub11_result_r_w),
			.i_fld_u_0_addr_0 (w_sub11_u_addr),
			.i_fld_u_0_datain_0 (w_sub11_u_datain),
			.o_fld_u_0_dataout_0 (w_sub11_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub11_u_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_result_1_addr_0 (w_sub14_result_addr),
			.i_fld_result_1_datain_0 (w_sub14_result_datain),
			.o_fld_result_1_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub14_result_r_w),
			.i_fld_u_0_addr_0 (w_sub14_u_addr),
			.i_fld_u_0_datain_0 (w_sub14_u_datain),
			.o_fld_u_0_dataout_0 (w_sub14_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub14_u_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_result_1_addr_0 (w_sub13_result_addr),
			.i_fld_result_1_datain_0 (w_sub13_result_datain),
			.o_fld_result_1_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub13_result_r_w),
			.i_fld_u_0_addr_0 (w_sub13_u_addr),
			.i_fld_u_0_datain_0 (w_sub13_u_datain),
			.o_fld_u_0_dataout_0 (w_sub13_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub13_u_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_result_1_addr_0 (w_sub15_result_addr),
			.i_fld_result_1_datain_0 (w_sub15_result_datain),
			.o_fld_result_1_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub15_result_r_w),
			.i_fld_u_0_addr_0 (w_sub15_u_addr),
			.i_fld_u_0_datain_0 (w_sub15_u_datain),
			.o_fld_u_0_dataout_0 (w_sub15_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub15_u_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_result_1_addr_0 (w_sub05_result_addr),
			.i_fld_result_1_datain_0 (w_sub05_result_datain),
			.o_fld_result_1_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_result_1_addr_0 (w_sub10_result_addr),
			.i_fld_result_1_datain_0 (w_sub10_result_datain),
			.o_fld_result_1_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub10_result_r_w),
			.i_fld_u_0_addr_0 (w_sub10_u_addr),
			.i_fld_u_0_datain_0 (w_sub10_u_datain),
			.o_fld_u_0_dataout_0 (w_sub10_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub10_u_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(10), .WORDS(1024) )
		dpram_uu_1(
			.clk (clock),
			.ce_0 (w_fld_uu_1_ce_0),
			.addr_0 (w_fld_uu_1_addr_0),
			.datain_0 (w_fld_uu_1_datain_0),
			.dataout_0 (w_fld_uu_1_dataout_0),
			.r_w_0 (w_fld_uu_1_r_w_0),
			.ce_1 (w_fld_uu_1_ce_1),
			.addr_1 (r_fld_uu_1_addr_1),
			.datain_1 (r_fld_uu_1_datain_1),
			.dataout_1 (w_fld_uu_1_dataout_1),
			.r_w_1 (r_fld_uu_1_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h35: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp94) ? 6'h14 : 6'h35);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp97) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1b)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp261) ? 6'h1e : 6'h20);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h34)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp573) ? 6'h24 : 6'h25);

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 6'h27;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 6'h29;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp681) ? 6'h2d : 6'h2f);

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1c)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp824) ? 6'h33 : 6'h11);

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h35: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h34)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1c)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1b)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h34)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h33)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h11)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1c)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1b)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h9)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h35: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp11[9:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp101[9:0] );

									end
									else
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp105[9:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp115[9:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp110[9:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp464[9:0] );

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp362[9:0] );

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp374[9:0] );

									end
									else
									if((r_sys_run_step==6'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp452[9:0] );

									end
									else
									if((r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp536[9:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp332[9:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp278[9:0] );

									end
									else
									if((r_sys_run_step==6'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp476[9:0] );

									end
									else
									if((r_sys_run_step==6'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp554[9:0] );

									end
									else
									if((r_sys_run_step==6'h28) || (r_sys_run_step==6'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp506[9:0] );

									end
									else
									if((r_sys_run_step==6'h29) || (r_sys_run_step==6'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp512[9:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp308[9:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp350[9:0] );

									end
									else
									if((r_sys_run_step==6'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp560[9:0] );

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp368[9:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp302[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp266[9:0] );

									end
									else
									if((r_sys_run_step==6'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp458[9:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp326[9:0] );

									end
									else
									if((r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp428[9:0] );

									end
									else
									if((r_sys_run_step==6'h14) || (r_sys_run_step==6'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp386[9:0] );

									end
									else
									if((r_sys_run_step==6'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp566[9:0] );

									end
									else
									if((r_sys_run_step==6'h17) || (r_sys_run_step==6'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp404[9:0] );

									end
									else
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp410[9:0] );

									end
									else
									if((r_sys_run_step==6'h25) || (r_sys_run_step==6'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp488[9:0] );

									end
									else
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp380[9:0] );

									end
									else
									if((r_sys_run_step==6'h24) || (r_sys_run_step==6'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp482[9:0] );

									end
									else
									if((r_sys_run_step==6'h1c) || (r_sys_run_step==6'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp434[9:0] );

									end
									else
									if((r_sys_run_step==6'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp470[9:0] );

									end
									else
									if((r_sys_run_step==6'h2c) || (r_sys_run_step==6'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp530[9:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp356[9:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp284[9:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp272[9:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp620[9:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp584[9:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp596[9:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp668[9:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp662[9:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp614[9:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp590[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp578[9:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp644[9:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp638[9:0] );

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp674[9:0] );

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp763[9:0] );

									end
									else
									if((r_sys_run_step==6'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp798[9:0] );

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp803[9:0] );

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp768[9:0] );

									end
									else
									if((r_sys_run_step==6'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp698[9:0] );

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp738[9:0] );

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp808[9:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp692[9:0] );

									end
									else
									if((r_sys_run_step==6'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp778[9:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp748[9:0] );

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp718[9:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp733[9:0] );

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp758[9:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp713[9:0] );

									end
									else
									if((r_sys_run_step==6'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp818[9:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp708[9:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp686[9:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp793[9:0] );

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp788[9:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp773[9:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp753[9:0] );

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp783[9:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp728[9:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp723[9:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp743[9:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp703[9:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp813[9:0] );

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp861[9:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp866[9:0] );

									end
									else
									if((r_sys_run_step==6'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp841[9:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp871[9:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp856[9:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp851[9:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp846[9:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp835[9:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp829[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp14;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp103;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp113;

									end
									else
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp108;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'ha)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==6'h14)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==6'h18)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h3)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp688;

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h1c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h3)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp831;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h32)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h10)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'ha)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h35: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_addr_1 <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp16[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_uu_1_datain_1 <= w_sys_tmp14;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h35: begin
							r_fld_uu_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_18 <= w_sys_tmp6;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_18 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h34)) begin
										r_run_k_18 <= w_sys_tmp571;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_18 <= w_sys_tmp572;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_run_k_18 <= w_sys_tmp679;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_18 <= w_sys_tmp680;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1c)) begin
										r_run_k_18 <= w_sys_tmp822;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_18 <= w_sys_tmp823;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_run_k_18 <= w_sys_tmp875;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_19 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_19 <= w_sys_tmp21;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_19 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h18)) begin
										r_run_j_19 <= w_sys_tmp122;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_20 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_20 <= w_sys_tmp96;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_mx_21 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_my_22 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_nlast_23 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_24 <= r_run_j_19;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_24 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_25 <= r_run_j_19;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1b)) begin
										r_run_copy0_j_25 <= w_sys_tmp119;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_26 <= r_run_j_19;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1a)) begin
										r_run_copy1_j_26 <= w_sys_tmp120;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_27 <= r_run_j_19;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h19)) begin
										r_run_copy2_j_27 <= w_sys_tmp121;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp488[9:0] );

									end
									else
									if((r_sys_run_step==6'h28)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp482[9:0] );

									end
									else
									if((r_sys_run_step==6'h2a)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp506[9:0] );

									end
									else
									if((r_sys_run_step==6'h2b)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp512[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h28<=r_sys_run_step && r_sys_run_step<=6'h2b)) begin
										r_sub09_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h28<=r_sys_run_step && r_sys_run_step<=6'h2b)) begin
										r_sub09_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub09_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp788[9:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp793[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h27)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp488[9:0] );

									end
									else
									if((r_sys_run_step==6'h25)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp476[9:0] );

									end
									else
									if((r_sys_run_step==6'h26)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp482[9:0] );

									end
									else
									if((r_sys_run_step==6'h24)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp470[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h24<=r_sys_run_step && r_sys_run_step<=6'h27)) begin
										r_sub08_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h24<=r_sys_run_step && r_sys_run_step<=6'h27)) begin
										r_sub08_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub08_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp783[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp778[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp584[9:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp596[9:0] );

									end
									else
									if((r_sys_run_step==6'h4)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp590[9:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp578[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sub12_u_datain <= w_sys_tmp580;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sub12_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub12_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp835[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp829[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp362[9:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp326[9:0] );

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp350[9:0] );

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp356[9:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp332[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'he<=r_sys_run_step && r_sys_run_step<=6'h12)) begin
										r_sub03_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'he<=r_sys_run_step && r_sys_run_step<=6'h12)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp728[9:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp723[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp718[9:0] );

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp871[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp302[9:0] );

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp326[9:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp308[9:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp332[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'ha<=r_sys_run_step && r_sys_run_step<=6'hd)) begin
										r_sub02_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'ha<=r_sys_run_step && r_sys_run_step<=6'hd)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp713[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp708[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h32)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp554[9:0] );

									end
									else
									if((r_sys_run_step==6'h31)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp536[9:0] );

									end
									else
									if((r_sys_run_step==6'h30)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp530[9:0] );

									end
									else
									if((r_sys_run_step==6'h34)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp566[9:0] );

									end
									else
									if((r_sys_run_step==6'h33)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp560[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h30<=r_sys_run_step && r_sys_run_step<=6'h34)) begin
										r_sub11_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h30<=r_sys_run_step && r_sys_run_step<=6'h34)) begin
										r_sub11_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub11_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp818[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp808[9:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp813[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp620[9:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp614[9:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp644[9:0] );

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp638[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'ha<=r_sys_run_step && r_sys_run_step<=6'hd)) begin
										r_sub14_u_datain <= w_sys_tmp580;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'ha<=r_sys_run_step && r_sys_run_step<=6'hd)) begin
										r_sub14_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub14_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp856[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp851[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp302[9:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp308[9:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp284[9:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp278[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h6<=r_sys_run_step && r_sys_run_step<=6'h9)) begin
										r_sub01_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h6<=r_sys_run_step && r_sys_run_step<=6'h9)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp703[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp698[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp620[9:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp596[9:0] );

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp614[9:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp590[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h6<=r_sys_run_step && r_sys_run_step<=6'h9)) begin
										r_sub13_u_datain <= w_sys_tmp580;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h6<=r_sys_run_step && r_sys_run_step<=6'h9)) begin
										r_sub13_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub13_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp841[9:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp846[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp266[9:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp284[9:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp272[9:0] );

									end
									else
									if((r_sys_run_step==6'h4)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp278[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sub00_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp692[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp686[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h23)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp464[9:0] );

									end
									else
									if((r_sys_run_step==6'h22)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp458[9:0] );

									end
									else
									if((r_sys_run_step==6'h20)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp434[9:0] );

									end
									else
									if((r_sys_run_step==6'h21)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp452[9:0] );

									end
									else
									if((r_sys_run_step==6'h1f)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp428[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h1f<=r_sys_run_step && r_sys_run_step<=6'h23)) begin
										r_sub07_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h1f<=r_sys_run_step && r_sys_run_step<=6'h23)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp763[9:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp773[9:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp768[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1c)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp410[9:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp404[9:0] );

									end
									else
									if((r_sys_run_step==6'h1e)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp434[9:0] );

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp428[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h1b<=r_sys_run_step && r_sys_run_step<=6'h1e)) begin
										r_sub06_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h1b<=r_sys_run_step && r_sys_run_step<=6'h1e)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp753[9:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp758[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp668[9:0] );

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp662[9:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp644[9:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp638[9:0] );

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp674[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'he<=r_sys_run_step && r_sys_run_step<=6'h12)) begin
										r_sub15_u_datain <= w_sys_tmp580;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'he<=r_sys_run_step && r_sys_run_step<=6'h12)) begin
										r_sub15_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub15_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp861[9:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp866[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp410[9:0] );

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp404[9:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp380[9:0] );

									end
									else
									if((r_sys_run_step==6'h18)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp386[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h17<=r_sys_run_step && r_sys_run_step<=6'h1a)) begin
										r_sub05_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h17<=r_sys_run_step && r_sys_run_step<=6'h1a)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp748[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp743[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h14)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp374[9:0] );

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp380[9:0] );

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp386[9:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp368[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h13<=r_sys_run_step && r_sys_run_step<=6'h16)) begin
										r_sub04_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h13<=r_sys_run_step && r_sys_run_step<=6'h16)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp733[9:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp738[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2f)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp536[9:0] );

									end
									else
									if((r_sys_run_step==6'h2c)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp506[9:0] );

									end
									else
									if((r_sys_run_step==6'h2d)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp512[9:0] );

									end
									else
									if((r_sys_run_step==6'h2e)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp530[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2c<=r_sys_run_step && r_sys_run_step<=6'h2f)) begin
										r_sub10_u_datain <= w_sys_tmp268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2c<=r_sys_run_step && r_sys_run_step<=6'h2f)) begin
										r_sub10_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub10_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp803[9:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp798[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h35: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp0_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp0_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp1_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp1_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp2_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp2_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp3_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp4_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp5_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp6_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp6_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp7_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp8_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp9_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp10_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp11_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp12_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp13_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp14_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp15_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp16_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp17_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp18_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp19_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp20_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp21_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp22_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp23_float <= w_sub03_result_dataout;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp23_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
