/*
TimeStamp:	2016/10/17		12:54
*/


module P3_2dim(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 3:0] r_sys_run_stage;
	reg         [ 5:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 3:0] w_sys_run_stage_p1;
	wire        [ 5:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [14:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [14:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [14:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [14:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [14:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [14:0] w_fld_V_3_addr_0;
	wire        [31:0] w_fld_V_3_datain_0;
	wire        [31:0] w_fld_V_3_dataout_0;
	wire               w_fld_V_3_r_w_0;
	wire               w_fld_V_3_ce_0;
	reg  signed [14:0] r_fld_V_3_addr_1;
	reg         [31:0] r_fld_V_3_datain_1;
	wire        [31:0] w_fld_V_3_dataout_1;
	reg                r_fld_V_3_r_w_1;
	wire               w_fld_V_3_ce_1;
	reg  signed [31:0] r_run_k_12;
	reg  signed [31:0] r_run_j_13;
	reg  signed [31:0] r_run_n_14;
	reg  signed [31:0] r_run_mx_15;
	reg  signed [31:0] r_run_my_16;
	reg         [31:0] r_run_dt_17;
	reg         [31:0] r_run_dx_18;
	reg         [31:0] r_run_dy_19;
	reg         [31:0] r_run_r1_20;
	reg         [31:0] r_run_r2_21;
	reg         [31:0] r_run_r3_22;
	reg         [31:0] r_run_r4_23;
	reg         [31:0] r_run_YY_24;
	reg  signed [31:0] r_run_kx_25;
	reg  signed [31:0] r_run_ky_26;
	reg  signed [31:0] r_run_nlast_27;
	reg  signed [31:0] r_run_copy0_j_28;
	reg  signed [31:0] r_run_copy1_j_29;
	reg  signed [31:0] r_run_copy2_j_30;
	reg  signed [31:0] r_run_copy0_j_31;
	reg  signed [31:0] r_run_copy1_j_32;
	reg  signed [31:0] r_run_copy2_j_33;
	reg  signed [31:0] r_run_copy3_j_34;
	reg  signed [31:0] r_run_copy4_j_35;
	reg  signed [31:0] r_run_copy0_j_36;
	reg  signed [31:0] r_run_copy1_j_37;
	reg  signed [31:0] r_run_copy2_j_38;
	reg  signed [31:0] r_run_copy3_j_39;
	reg  signed [31:0] r_run_copy4_j_40;
	reg  signed [31:0] r_run_copy0_j_41;
	reg  signed [31:0] r_run_copy1_j_42;
	reg  signed [31:0] r_run_copy2_j_43;
	reg  signed [31:0] r_run_copy3_j_44;
	reg  signed [31:0] r_run_copy4_j_45;
	reg  signed [31:0] r_run_copy0_j_46;
	reg  signed [31:0] r_run_copy1_j_47;
	reg  signed [31:0] r_run_copy2_j_48;
	reg  signed [31:0] r_run_copy3_j_49;
	reg  signed [31:0] r_run_copy4_j_50;
	reg  signed [31:0] r_run_copy0_j_51;
	reg  signed [31:0] r_run_copy1_j_52;
	reg  signed [31:0] r_run_copy2_j_53;
	reg  signed [31:0] r_run_copy3_j_54;
	reg  signed [31:0] r_run_copy4_j_55;
	reg  signed [31:0] r_run_copy0_j_56;
	reg  signed [31:0] r_run_copy1_j_57;
	reg  signed [31:0] r_run_copy2_j_58;
	reg  signed [31:0] r_run_copy3_j_59;
	reg  signed [31:0] r_run_copy4_j_60;
	reg  signed [31:0] r_run_copy0_j_61;
	reg  signed [31:0] r_run_copy1_j_62;
	reg  signed [31:0] r_run_copy2_j_63;
	reg  signed [31:0] r_run_copy3_j_64;
	reg  signed [31:0] r_run_copy4_j_65;
	reg  signed [31:0] r_run_copy0_j_66;
	reg  signed [31:0] r_run_copy1_j_67;
	reg  signed [31:0] r_run_copy2_j_68;
	reg  signed [31:0] r_run_copy3_j_69;
	reg  signed [31:0] r_run_copy4_j_70;
	reg  signed [31:0] r_run_copy0_j_71;
	reg  signed [31:0] r_run_copy1_j_72;
	reg  signed [31:0] r_run_copy2_j_73;
	reg  signed [31:0] r_run_copy0_j_74;
	reg  signed [31:0] r_run_copy1_j_75;
	reg  signed [31:0] r_run_copy2_j_76;
	reg  signed [31:0] r_run_copy0_j_77;
	reg  signed [31:0] r_run_copy1_j_78;
	reg  signed [31:0] r_run_copy2_j_79;
	reg  signed [31:0] r_run_copy0_j_80;
	reg  signed [31:0] r_run_copy1_j_81;
	reg  signed [31:0] r_run_copy2_j_82;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 8:0] w_sub03_T_addr;
	reg  signed [ 8:0] r_sub03_T_addr;
	wire        [31:0] w_sub03_T_datain;
	reg         [31:0] r_sub03_T_datain;
	wire        [31:0] w_sub03_T_dataout;
	wire               w_sub03_T_r_w;
	reg                r_sub03_T_r_w;
	wire signed [ 8:0] w_sub03_V_addr;
	reg  signed [ 8:0] r_sub03_V_addr;
	wire        [31:0] w_sub03_V_datain;
	reg         [31:0] r_sub03_V_datain;
	wire        [31:0] w_sub03_V_dataout;
	wire               w_sub03_V_r_w;
	reg                r_sub03_V_r_w;
	wire signed [ 8:0] w_sub03_U_addr;
	reg  signed [ 8:0] r_sub03_U_addr;
	wire        [31:0] w_sub03_U_datain;
	reg         [31:0] r_sub03_U_datain;
	wire        [31:0] w_sub03_U_dataout;
	wire               w_sub03_U_r_w;
	reg                r_sub03_U_r_w;
	wire signed [ 8:0] w_sub03_result_addr;
	reg  signed [ 8:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 8:0] w_sub02_T_addr;
	reg  signed [ 8:0] r_sub02_T_addr;
	wire        [31:0] w_sub02_T_datain;
	reg         [31:0] r_sub02_T_datain;
	wire        [31:0] w_sub02_T_dataout;
	wire               w_sub02_T_r_w;
	reg                r_sub02_T_r_w;
	wire signed [ 8:0] w_sub02_V_addr;
	reg  signed [ 8:0] r_sub02_V_addr;
	wire        [31:0] w_sub02_V_datain;
	reg         [31:0] r_sub02_V_datain;
	wire        [31:0] w_sub02_V_dataout;
	wire               w_sub02_V_r_w;
	reg                r_sub02_V_r_w;
	wire signed [ 8:0] w_sub02_U_addr;
	reg  signed [ 8:0] r_sub02_U_addr;
	wire        [31:0] w_sub02_U_datain;
	reg         [31:0] r_sub02_U_datain;
	wire        [31:0] w_sub02_U_dataout;
	wire               w_sub02_U_r_w;
	reg                r_sub02_U_r_w;
	wire signed [ 8:0] w_sub02_result_addr;
	reg  signed [ 8:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 8:0] w_sub01_T_addr;
	reg  signed [ 8:0] r_sub01_T_addr;
	wire        [31:0] w_sub01_T_datain;
	reg         [31:0] r_sub01_T_datain;
	wire        [31:0] w_sub01_T_dataout;
	wire               w_sub01_T_r_w;
	reg                r_sub01_T_r_w;
	wire signed [ 8:0] w_sub01_V_addr;
	reg  signed [ 8:0] r_sub01_V_addr;
	wire        [31:0] w_sub01_V_datain;
	reg         [31:0] r_sub01_V_datain;
	wire        [31:0] w_sub01_V_dataout;
	wire               w_sub01_V_r_w;
	reg                r_sub01_V_r_w;
	wire signed [ 8:0] w_sub01_U_addr;
	reg  signed [ 8:0] r_sub01_U_addr;
	wire        [31:0] w_sub01_U_datain;
	reg         [31:0] r_sub01_U_datain;
	wire        [31:0] w_sub01_U_dataout;
	wire               w_sub01_U_r_w;
	reg                r_sub01_U_r_w;
	wire signed [ 8:0] w_sub01_result_addr;
	reg  signed [ 8:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [14:0] w_sub00_T_addr;
	reg  signed [14:0] r_sub00_T_addr;
	wire        [31:0] w_sub00_T_datain;
	reg         [31:0] r_sub00_T_datain;
	wire        [31:0] w_sub00_T_dataout;
	wire               w_sub00_T_r_w;
	reg                r_sub00_T_r_w;
	wire signed [14:0] w_sub00_V_addr;
	reg  signed [14:0] r_sub00_V_addr;
	wire        [31:0] w_sub00_V_datain;
	reg         [31:0] r_sub00_V_datain;
	wire        [31:0] w_sub00_V_dataout;
	wire               w_sub00_V_r_w;
	reg                r_sub00_V_r_w;
	wire signed [14:0] w_sub00_U_addr;
	reg  signed [14:0] r_sub00_U_addr;
	wire        [31:0] w_sub00_U_datain;
	reg         [31:0] r_sub00_U_datain;
	wire        [31:0] w_sub00_U_dataout;
	wire               w_sub00_U_r_w;
	reg                r_sub00_U_r_w;
	wire signed [14:0] w_sub00_result_addr;
	reg  signed [14:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [ 8:0] w_sub07_T_addr;
	reg  signed [ 8:0] r_sub07_T_addr;
	wire        [31:0] w_sub07_T_datain;
	reg         [31:0] r_sub07_T_datain;
	wire        [31:0] w_sub07_T_dataout;
	wire               w_sub07_T_r_w;
	reg                r_sub07_T_r_w;
	wire signed [ 8:0] w_sub07_V_addr;
	reg  signed [ 8:0] r_sub07_V_addr;
	wire        [31:0] w_sub07_V_datain;
	reg         [31:0] r_sub07_V_datain;
	wire        [31:0] w_sub07_V_dataout;
	wire               w_sub07_V_r_w;
	reg                r_sub07_V_r_w;
	wire signed [ 8:0] w_sub07_U_addr;
	reg  signed [ 8:0] r_sub07_U_addr;
	wire        [31:0] w_sub07_U_datain;
	reg         [31:0] r_sub07_U_datain;
	wire        [31:0] w_sub07_U_dataout;
	wire               w_sub07_U_r_w;
	reg                r_sub07_U_r_w;
	wire signed [ 8:0] w_sub07_result_addr;
	reg  signed [ 8:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [ 8:0] w_sub06_T_addr;
	reg  signed [ 8:0] r_sub06_T_addr;
	wire        [31:0] w_sub06_T_datain;
	reg         [31:0] r_sub06_T_datain;
	wire        [31:0] w_sub06_T_dataout;
	wire               w_sub06_T_r_w;
	reg                r_sub06_T_r_w;
	wire signed [ 8:0] w_sub06_V_addr;
	reg  signed [ 8:0] r_sub06_V_addr;
	wire        [31:0] w_sub06_V_datain;
	reg         [31:0] r_sub06_V_datain;
	wire        [31:0] w_sub06_V_dataout;
	wire               w_sub06_V_r_w;
	reg                r_sub06_V_r_w;
	wire signed [ 8:0] w_sub06_U_addr;
	reg  signed [ 8:0] r_sub06_U_addr;
	wire        [31:0] w_sub06_U_datain;
	reg         [31:0] r_sub06_U_datain;
	wire        [31:0] w_sub06_U_dataout;
	wire               w_sub06_U_r_w;
	reg                r_sub06_U_r_w;
	wire signed [ 8:0] w_sub06_result_addr;
	reg  signed [ 8:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [ 8:0] w_sub05_T_addr;
	reg  signed [ 8:0] r_sub05_T_addr;
	wire        [31:0] w_sub05_T_datain;
	reg         [31:0] r_sub05_T_datain;
	wire        [31:0] w_sub05_T_dataout;
	wire               w_sub05_T_r_w;
	reg                r_sub05_T_r_w;
	wire signed [ 8:0] w_sub05_V_addr;
	reg  signed [ 8:0] r_sub05_V_addr;
	wire        [31:0] w_sub05_V_datain;
	reg         [31:0] r_sub05_V_datain;
	wire        [31:0] w_sub05_V_dataout;
	wire               w_sub05_V_r_w;
	reg                r_sub05_V_r_w;
	wire signed [ 8:0] w_sub05_U_addr;
	reg  signed [ 8:0] r_sub05_U_addr;
	wire        [31:0] w_sub05_U_datain;
	reg         [31:0] r_sub05_U_datain;
	wire        [31:0] w_sub05_U_dataout;
	wire               w_sub05_U_r_w;
	reg                r_sub05_U_r_w;
	wire signed [ 8:0] w_sub05_result_addr;
	reg  signed [ 8:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [ 8:0] w_sub04_T_addr;
	reg  signed [ 8:0] r_sub04_T_addr;
	wire        [31:0] w_sub04_T_datain;
	reg         [31:0] r_sub04_T_datain;
	wire        [31:0] w_sub04_T_dataout;
	wire               w_sub04_T_r_w;
	reg                r_sub04_T_r_w;
	wire signed [ 8:0] w_sub04_V_addr;
	reg  signed [ 8:0] r_sub04_V_addr;
	wire        [31:0] w_sub04_V_datain;
	reg         [31:0] r_sub04_V_datain;
	wire        [31:0] w_sub04_V_dataout;
	wire               w_sub04_V_r_w;
	reg                r_sub04_V_r_w;
	wire signed [ 8:0] w_sub04_U_addr;
	reg  signed [ 8:0] r_sub04_U_addr;
	wire        [31:0] w_sub04_U_datain;
	reg         [31:0] r_sub04_U_datain;
	wire        [31:0] w_sub04_U_dataout;
	wire               w_sub04_U_r_w;
	reg                r_sub04_U_r_w;
	wire signed [ 8:0] w_sub04_result_addr;
	reg  signed [ 8:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire               w_sys_tmp12;
	wire               w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp15;
	wire               w_sys_tmp16;
	wire        [31:0] w_sys_tmp18;
	wire        [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire        [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp27;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp32;
	wire signed [31:0] w_sys_tmp33;
	wire        [31:0] w_sys_tmp36;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp45;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire        [31:0] w_sys_tmp128;
	wire               w_sys_tmp226;
	wire               w_sys_tmp227;
	wire signed [31:0] w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire               w_sys_tmp230;
	wire               w_sys_tmp231;
	wire signed [31:0] w_sys_tmp232;
	wire signed [31:0] w_sys_tmp235;
	wire signed [31:0] w_sys_tmp236;
	wire signed [31:0] w_sys_tmp237;
	wire        [31:0] w_sys_tmp238;
	wire signed [31:0] w_sys_tmp239;
	wire signed [31:0] w_sys_tmp240;
	wire signed [31:0] w_sys_tmp243;
	wire signed [31:0] w_sys_tmp244;
	wire        [31:0] w_sys_tmp246;
	wire signed [31:0] w_sys_tmp247;
	wire signed [31:0] w_sys_tmp248;
	wire signed [31:0] w_sys_tmp251;
	wire signed [31:0] w_sys_tmp252;
	wire        [31:0] w_sys_tmp254;
	wire signed [31:0] w_sys_tmp255;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp258;
	wire signed [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp260;
	wire signed [31:0] w_sys_tmp261;
	wire signed [31:0] w_sys_tmp262;
	wire signed [31:0] w_sys_tmp263;
	wire signed [31:0] w_sys_tmp444;
	wire               w_sys_tmp445;
	wire               w_sys_tmp446;
	wire signed [31:0] w_sys_tmp447;
	wire signed [31:0] w_sys_tmp450;
	wire signed [31:0] w_sys_tmp451;
	wire signed [31:0] w_sys_tmp452;
	wire        [31:0] w_sys_tmp453;
	wire signed [31:0] w_sys_tmp454;
	wire signed [31:0] w_sys_tmp455;
	wire signed [31:0] w_sys_tmp458;
	wire signed [31:0] w_sys_tmp459;
	wire        [31:0] w_sys_tmp461;
	wire signed [31:0] w_sys_tmp462;
	wire signed [31:0] w_sys_tmp463;
	wire signed [31:0] w_sys_tmp466;
	wire signed [31:0] w_sys_tmp467;
	wire        [31:0] w_sys_tmp469;
	wire signed [31:0] w_sys_tmp470;
	wire signed [31:0] w_sys_tmp471;
	wire signed [31:0] w_sys_tmp473;
	wire signed [31:0] w_sys_tmp474;
	wire signed [31:0] w_sys_tmp475;
	wire signed [31:0] w_sys_tmp476;
	wire signed [31:0] w_sys_tmp477;
	wire signed [31:0] w_sys_tmp478;
	wire signed [31:0] w_sys_tmp659;
	wire               w_sys_tmp660;
	wire               w_sys_tmp661;
	wire signed [31:0] w_sys_tmp662;
	wire signed [31:0] w_sys_tmp665;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp667;
	wire        [31:0] w_sys_tmp668;
	wire signed [31:0] w_sys_tmp669;
	wire signed [31:0] w_sys_tmp670;
	wire signed [31:0] w_sys_tmp673;
	wire signed [31:0] w_sys_tmp674;
	wire        [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp677;
	wire signed [31:0] w_sys_tmp678;
	wire signed [31:0] w_sys_tmp681;
	wire signed [31:0] w_sys_tmp682;
	wire        [31:0] w_sys_tmp684;
	wire signed [31:0] w_sys_tmp685;
	wire signed [31:0] w_sys_tmp686;
	wire signed [31:0] w_sys_tmp688;
	wire signed [31:0] w_sys_tmp689;
	wire signed [31:0] w_sys_tmp690;
	wire signed [31:0] w_sys_tmp691;
	wire signed [31:0] w_sys_tmp692;
	wire signed [31:0] w_sys_tmp693;
	wire signed [31:0] w_sys_tmp874;
	wire               w_sys_tmp875;
	wire               w_sys_tmp876;
	wire signed [31:0] w_sys_tmp877;
	wire signed [31:0] w_sys_tmp880;
	wire signed [31:0] w_sys_tmp881;
	wire signed [31:0] w_sys_tmp882;
	wire        [31:0] w_sys_tmp883;
	wire signed [31:0] w_sys_tmp884;
	wire signed [31:0] w_sys_tmp885;
	wire signed [31:0] w_sys_tmp888;
	wire signed [31:0] w_sys_tmp889;
	wire        [31:0] w_sys_tmp891;
	wire signed [31:0] w_sys_tmp892;
	wire signed [31:0] w_sys_tmp893;
	wire signed [31:0] w_sys_tmp896;
	wire signed [31:0] w_sys_tmp897;
	wire        [31:0] w_sys_tmp899;
	wire signed [31:0] w_sys_tmp900;
	wire signed [31:0] w_sys_tmp901;
	wire signed [31:0] w_sys_tmp903;
	wire signed [31:0] w_sys_tmp904;
	wire signed [31:0] w_sys_tmp905;
	wire signed [31:0] w_sys_tmp906;
	wire signed [31:0] w_sys_tmp907;
	wire signed [31:0] w_sys_tmp908;
	wire signed [31:0] w_sys_tmp1089;
	wire               w_sys_tmp1090;
	wire               w_sys_tmp1091;
	wire signed [31:0] w_sys_tmp1092;
	wire signed [31:0] w_sys_tmp1093;
	wire               w_sys_tmp1094;
	wire               w_sys_tmp1095;
	wire signed [31:0] w_sys_tmp1096;
	wire signed [31:0] w_sys_tmp1099;
	wire signed [31:0] w_sys_tmp1100;
	wire signed [31:0] w_sys_tmp1101;
	wire        [31:0] w_sys_tmp1102;
	wire signed [31:0] w_sys_tmp1103;
	wire signed [31:0] w_sys_tmp1104;
	wire signed [31:0] w_sys_tmp1107;
	wire signed [31:0] w_sys_tmp1108;
	wire        [31:0] w_sys_tmp1110;
	wire signed [31:0] w_sys_tmp1111;
	wire signed [31:0] w_sys_tmp1112;
	wire signed [31:0] w_sys_tmp1115;
	wire signed [31:0] w_sys_tmp1116;
	wire        [31:0] w_sys_tmp1118;
	wire signed [31:0] w_sys_tmp1119;
	wire signed [31:0] w_sys_tmp1120;
	wire signed [31:0] w_sys_tmp1122;
	wire signed [31:0] w_sys_tmp1123;
	wire signed [31:0] w_sys_tmp1124;
	wire signed [31:0] w_sys_tmp1125;
	wire signed [31:0] w_sys_tmp1126;
	wire signed [31:0] w_sys_tmp1127;
	wire signed [31:0] w_sys_tmp1308;
	wire               w_sys_tmp1309;
	wire               w_sys_tmp1310;
	wire signed [31:0] w_sys_tmp1311;
	wire signed [31:0] w_sys_tmp1314;
	wire signed [31:0] w_sys_tmp1315;
	wire signed [31:0] w_sys_tmp1316;
	wire        [31:0] w_sys_tmp1317;
	wire signed [31:0] w_sys_tmp1318;
	wire signed [31:0] w_sys_tmp1319;
	wire signed [31:0] w_sys_tmp1322;
	wire signed [31:0] w_sys_tmp1323;
	wire        [31:0] w_sys_tmp1325;
	wire signed [31:0] w_sys_tmp1326;
	wire signed [31:0] w_sys_tmp1327;
	wire signed [31:0] w_sys_tmp1330;
	wire signed [31:0] w_sys_tmp1331;
	wire        [31:0] w_sys_tmp1333;
	wire signed [31:0] w_sys_tmp1334;
	wire signed [31:0] w_sys_tmp1335;
	wire signed [31:0] w_sys_tmp1337;
	wire signed [31:0] w_sys_tmp1338;
	wire signed [31:0] w_sys_tmp1339;
	wire signed [31:0] w_sys_tmp1340;
	wire signed [31:0] w_sys_tmp1341;
	wire signed [31:0] w_sys_tmp1342;
	wire signed [31:0] w_sys_tmp1523;
	wire               w_sys_tmp1524;
	wire               w_sys_tmp1525;
	wire signed [31:0] w_sys_tmp1526;
	wire signed [31:0] w_sys_tmp1529;
	wire signed [31:0] w_sys_tmp1530;
	wire signed [31:0] w_sys_tmp1531;
	wire        [31:0] w_sys_tmp1532;
	wire signed [31:0] w_sys_tmp1533;
	wire signed [31:0] w_sys_tmp1534;
	wire signed [31:0] w_sys_tmp1537;
	wire signed [31:0] w_sys_tmp1538;
	wire        [31:0] w_sys_tmp1540;
	wire signed [31:0] w_sys_tmp1541;
	wire signed [31:0] w_sys_tmp1542;
	wire signed [31:0] w_sys_tmp1545;
	wire signed [31:0] w_sys_tmp1546;
	wire        [31:0] w_sys_tmp1548;
	wire signed [31:0] w_sys_tmp1549;
	wire signed [31:0] w_sys_tmp1550;
	wire signed [31:0] w_sys_tmp1552;
	wire signed [31:0] w_sys_tmp1553;
	wire signed [31:0] w_sys_tmp1554;
	wire signed [31:0] w_sys_tmp1555;
	wire signed [31:0] w_sys_tmp1556;
	wire signed [31:0] w_sys_tmp1557;
	wire signed [31:0] w_sys_tmp1738;
	wire               w_sys_tmp1739;
	wire               w_sys_tmp1740;
	wire signed [31:0] w_sys_tmp1741;
	wire signed [31:0] w_sys_tmp1744;
	wire signed [31:0] w_sys_tmp1745;
	wire signed [31:0] w_sys_tmp1746;
	wire        [31:0] w_sys_tmp1747;
	wire signed [31:0] w_sys_tmp1748;
	wire signed [31:0] w_sys_tmp1749;
	wire signed [31:0] w_sys_tmp1752;
	wire signed [31:0] w_sys_tmp1753;
	wire        [31:0] w_sys_tmp1755;
	wire signed [31:0] w_sys_tmp1756;
	wire signed [31:0] w_sys_tmp1757;
	wire signed [31:0] w_sys_tmp1760;
	wire signed [31:0] w_sys_tmp1761;
	wire        [31:0] w_sys_tmp1763;
	wire signed [31:0] w_sys_tmp1764;
	wire signed [31:0] w_sys_tmp1765;
	wire signed [31:0] w_sys_tmp1767;
	wire signed [31:0] w_sys_tmp1768;
	wire signed [31:0] w_sys_tmp1769;
	wire signed [31:0] w_sys_tmp1770;
	wire signed [31:0] w_sys_tmp1771;
	wire signed [31:0] w_sys_tmp1772;
	wire               w_sys_tmp1953;
	wire               w_sys_tmp1954;
	wire signed [31:0] w_sys_tmp1955;
	wire signed [31:0] w_sys_tmp1956;
	wire               w_sys_tmp1957;
	wire               w_sys_tmp1958;
	wire signed [31:0] w_sys_tmp1959;
	wire signed [31:0] w_sys_tmp1962;
	wire signed [31:0] w_sys_tmp1963;
	wire        [31:0] w_sys_tmp1964;
	wire signed [31:0] w_sys_tmp1968;
	wire signed [31:0] w_sys_tmp1969;
	wire        [31:0] w_sys_tmp1970;
	wire signed [31:0] w_sys_tmp1974;
	wire signed [31:0] w_sys_tmp1975;
	wire        [31:0] w_sys_tmp1976;
	wire signed [31:0] w_sys_tmp1980;
	wire signed [31:0] w_sys_tmp1981;
	wire signed [31:0] w_sys_tmp1985;
	wire signed [31:0] w_sys_tmp1986;
	wire signed [31:0] w_sys_tmp1990;
	wire signed [31:0] w_sys_tmp1991;
	wire signed [31:0] w_sys_tmp1994;
	wire signed [31:0] w_sys_tmp1995;
	wire               w_sys_tmp1996;
	wire               w_sys_tmp1997;
	wire signed [31:0] w_sys_tmp1998;
	wire signed [31:0] w_sys_tmp2001;
	wire signed [31:0] w_sys_tmp2002;
	wire signed [31:0] w_sys_tmp2003;
	wire signed [31:0] w_sys_tmp2004;
	wire        [31:0] w_sys_tmp2005;
	wire signed [31:0] w_sys_tmp2006;
	wire signed [31:0] w_sys_tmp2007;
	wire signed [31:0] w_sys_tmp2011;
	wire signed [31:0] w_sys_tmp2012;
	wire signed [31:0] w_sys_tmp2014;
	wire        [31:0] w_sys_tmp2015;
	wire signed [31:0] w_sys_tmp2016;
	wire signed [31:0] w_sys_tmp2017;
	wire signed [31:0] w_sys_tmp2020;
	wire signed [31:0] w_sys_tmp2021;
	wire signed [31:0] w_sys_tmp2022;
	wire signed [31:0] w_sys_tmp2023;
	wire signed [31:0] w_sys_tmp2168;
	wire               w_sys_tmp2169;
	wire               w_sys_tmp2170;
	wire signed [31:0] w_sys_tmp2171;
	wire signed [31:0] w_sys_tmp2174;
	wire signed [31:0] w_sys_tmp2175;
	wire signed [31:0] w_sys_tmp2176;
	wire signed [31:0] w_sys_tmp2177;
	wire        [31:0] w_sys_tmp2178;
	wire signed [31:0] w_sys_tmp2179;
	wire signed [31:0] w_sys_tmp2180;
	wire signed [31:0] w_sys_tmp2184;
	wire signed [31:0] w_sys_tmp2185;
	wire signed [31:0] w_sys_tmp2187;
	wire        [31:0] w_sys_tmp2188;
	wire signed [31:0] w_sys_tmp2189;
	wire signed [31:0] w_sys_tmp2190;
	wire signed [31:0] w_sys_tmp2193;
	wire signed [31:0] w_sys_tmp2194;
	wire signed [31:0] w_sys_tmp2195;
	wire signed [31:0] w_sys_tmp2196;
	wire signed [31:0] w_sys_tmp2341;
	wire               w_sys_tmp2342;
	wire               w_sys_tmp2343;
	wire signed [31:0] w_sys_tmp2344;
	wire signed [31:0] w_sys_tmp2347;
	wire signed [31:0] w_sys_tmp2348;
	wire signed [31:0] w_sys_tmp2349;
	wire signed [31:0] w_sys_tmp2350;
	wire        [31:0] w_sys_tmp2351;
	wire signed [31:0] w_sys_tmp2352;
	wire signed [31:0] w_sys_tmp2353;
	wire signed [31:0] w_sys_tmp2357;
	wire signed [31:0] w_sys_tmp2358;
	wire signed [31:0] w_sys_tmp2360;
	wire        [31:0] w_sys_tmp2361;
	wire signed [31:0] w_sys_tmp2362;
	wire signed [31:0] w_sys_tmp2363;
	wire signed [31:0] w_sys_tmp2366;
	wire signed [31:0] w_sys_tmp2367;
	wire signed [31:0] w_sys_tmp2368;
	wire signed [31:0] w_sys_tmp2369;
	wire signed [31:0] w_sys_tmp2514;
	wire               w_sys_tmp2515;
	wire               w_sys_tmp2516;
	wire signed [31:0] w_sys_tmp2517;
	wire signed [31:0] w_sys_tmp2520;
	wire signed [31:0] w_sys_tmp2521;
	wire signed [31:0] w_sys_tmp2522;
	wire signed [31:0] w_sys_tmp2523;
	wire        [31:0] w_sys_tmp2524;
	wire signed [31:0] w_sys_tmp2525;
	wire signed [31:0] w_sys_tmp2526;
	wire signed [31:0] w_sys_tmp2530;
	wire signed [31:0] w_sys_tmp2531;
	wire signed [31:0] w_sys_tmp2533;
	wire        [31:0] w_sys_tmp2534;
	wire signed [31:0] w_sys_tmp2535;
	wire signed [31:0] w_sys_tmp2536;
	wire signed [31:0] w_sys_tmp2539;
	wire signed [31:0] w_sys_tmp2540;
	wire signed [31:0] w_sys_tmp2541;
	wire signed [31:0] w_sys_tmp2542;
	wire signed [31:0] w_sys_tmp2687;
	wire               w_sys_tmp2688;
	wire               w_sys_tmp2689;
	wire signed [31:0] w_sys_tmp2690;
	wire signed [31:0] w_sys_tmp2693;
	wire signed [31:0] w_sys_tmp2694;
	wire        [31:0] w_sys_tmp2695;
	wire signed [31:0] w_sys_tmp2699;
	wire signed [31:0] w_sys_tmp2700;
	wire        [31:0] w_sys_tmp2701;
	wire signed [31:0] w_sys_tmp2705;
	wire signed [31:0] w_sys_tmp2706;
	wire signed [31:0] w_sys_tmp2710;
	wire signed [31:0] w_sys_tmp2711;
	wire        [31:0] w_sys_tmp2712;
	wire signed [31:0] w_sys_tmp2716;
	wire signed [31:0] w_sys_tmp2717;
	wire signed [31:0] w_sys_tmp2722;
	wire signed [31:0] w_sys_tmp2723;
	wire signed [31:0] w_sys_tmp2726;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 4'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 6'h1);
	assign w_fld_T_0_addr_0 = 15'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 15'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 15'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_fld_V_3_addr_0 = 15'sh0;
	assign w_fld_V_3_datain_0 = 32'h0;
	assign w_fld_V_3_r_w_0 = 1'h0;
	assign w_fld_V_3_ce_0 = w_sys_ce;
	assign w_fld_V_3_ce_1 = w_sys_ce;
	assign w_sub03_T_addr = ( (|r_sys_processing_methodID) ? r_sub03_T_addr : 9'sh0 ) ;
	assign w_sub03_T_datain = ( (|r_sys_processing_methodID) ? r_sub03_T_datain : 32'h0 ) ;
	assign w_sub03_T_r_w = ( (|r_sys_processing_methodID) ? r_sub03_T_r_w : 1'h0 ) ;
	assign w_sub03_V_addr = ( (|r_sys_processing_methodID) ? r_sub03_V_addr : 9'sh0 ) ;
	assign w_sub03_V_datain = ( (|r_sys_processing_methodID) ? r_sub03_V_datain : 32'h0 ) ;
	assign w_sub03_V_r_w = ( (|r_sys_processing_methodID) ? r_sub03_V_r_w : 1'h0 ) ;
	assign w_sub03_U_addr = ( (|r_sys_processing_methodID) ? r_sub03_U_addr : 9'sh0 ) ;
	assign w_sub03_U_datain = ( (|r_sys_processing_methodID) ? r_sub03_U_datain : 32'h0 ) ;
	assign w_sub03_U_r_w = ( (|r_sys_processing_methodID) ? r_sub03_U_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 9'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_T_addr = ( (|r_sys_processing_methodID) ? r_sub02_T_addr : 9'sh0 ) ;
	assign w_sub02_T_datain = ( (|r_sys_processing_methodID) ? r_sub02_T_datain : 32'h0 ) ;
	assign w_sub02_T_r_w = ( (|r_sys_processing_methodID) ? r_sub02_T_r_w : 1'h0 ) ;
	assign w_sub02_V_addr = ( (|r_sys_processing_methodID) ? r_sub02_V_addr : 9'sh0 ) ;
	assign w_sub02_V_datain = ( (|r_sys_processing_methodID) ? r_sub02_V_datain : 32'h0 ) ;
	assign w_sub02_V_r_w = ( (|r_sys_processing_methodID) ? r_sub02_V_r_w : 1'h0 ) ;
	assign w_sub02_U_addr = ( (|r_sys_processing_methodID) ? r_sub02_U_addr : 9'sh0 ) ;
	assign w_sub02_U_datain = ( (|r_sys_processing_methodID) ? r_sub02_U_datain : 32'h0 ) ;
	assign w_sub02_U_r_w = ( (|r_sys_processing_methodID) ? r_sub02_U_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 9'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_T_addr = ( (|r_sys_processing_methodID) ? r_sub01_T_addr : 9'sh0 ) ;
	assign w_sub01_T_datain = ( (|r_sys_processing_methodID) ? r_sub01_T_datain : 32'h0 ) ;
	assign w_sub01_T_r_w = ( (|r_sys_processing_methodID) ? r_sub01_T_r_w : 1'h0 ) ;
	assign w_sub01_V_addr = ( (|r_sys_processing_methodID) ? r_sub01_V_addr : 9'sh0 ) ;
	assign w_sub01_V_datain = ( (|r_sys_processing_methodID) ? r_sub01_V_datain : 32'h0 ) ;
	assign w_sub01_V_r_w = ( (|r_sys_processing_methodID) ? r_sub01_V_r_w : 1'h0 ) ;
	assign w_sub01_U_addr = ( (|r_sys_processing_methodID) ? r_sub01_U_addr : 9'sh0 ) ;
	assign w_sub01_U_datain = ( (|r_sys_processing_methodID) ? r_sub01_U_datain : 32'h0 ) ;
	assign w_sub01_U_r_w = ( (|r_sys_processing_methodID) ? r_sub01_U_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 9'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_T_addr = ( (|r_sys_processing_methodID) ? r_sub00_T_addr : 15'sh0 ) ;
	assign w_sub00_T_datain = ( (|r_sys_processing_methodID) ? r_sub00_T_datain : 32'h0 ) ;
	assign w_sub00_T_r_w = ( (|r_sys_processing_methodID) ? r_sub00_T_r_w : 1'h0 ) ;
	assign w_sub00_V_addr = ( (|r_sys_processing_methodID) ? r_sub00_V_addr : 15'sh0 ) ;
	assign w_sub00_V_datain = ( (|r_sys_processing_methodID) ? r_sub00_V_datain : 32'h0 ) ;
	assign w_sub00_V_r_w = ( (|r_sys_processing_methodID) ? r_sub00_V_r_w : 1'h0 ) ;
	assign w_sub00_U_addr = ( (|r_sys_processing_methodID) ? r_sub00_U_addr : 15'sh0 ) ;
	assign w_sub00_U_datain = ( (|r_sys_processing_methodID) ? r_sub00_U_datain : 32'h0 ) ;
	assign w_sub00_U_r_w = ( (|r_sys_processing_methodID) ? r_sub00_U_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 15'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_T_addr = ( (|r_sys_processing_methodID) ? r_sub07_T_addr : 9'sh0 ) ;
	assign w_sub07_T_datain = ( (|r_sys_processing_methodID) ? r_sub07_T_datain : 32'h0 ) ;
	assign w_sub07_T_r_w = ( (|r_sys_processing_methodID) ? r_sub07_T_r_w : 1'h0 ) ;
	assign w_sub07_V_addr = ( (|r_sys_processing_methodID) ? r_sub07_V_addr : 9'sh0 ) ;
	assign w_sub07_V_datain = ( (|r_sys_processing_methodID) ? r_sub07_V_datain : 32'h0 ) ;
	assign w_sub07_V_r_w = ( (|r_sys_processing_methodID) ? r_sub07_V_r_w : 1'h0 ) ;
	assign w_sub07_U_addr = ( (|r_sys_processing_methodID) ? r_sub07_U_addr : 9'sh0 ) ;
	assign w_sub07_U_datain = ( (|r_sys_processing_methodID) ? r_sub07_U_datain : 32'h0 ) ;
	assign w_sub07_U_r_w = ( (|r_sys_processing_methodID) ? r_sub07_U_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 9'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_T_addr = ( (|r_sys_processing_methodID) ? r_sub06_T_addr : 9'sh0 ) ;
	assign w_sub06_T_datain = ( (|r_sys_processing_methodID) ? r_sub06_T_datain : 32'h0 ) ;
	assign w_sub06_T_r_w = ( (|r_sys_processing_methodID) ? r_sub06_T_r_w : 1'h0 ) ;
	assign w_sub06_V_addr = ( (|r_sys_processing_methodID) ? r_sub06_V_addr : 9'sh0 ) ;
	assign w_sub06_V_datain = ( (|r_sys_processing_methodID) ? r_sub06_V_datain : 32'h0 ) ;
	assign w_sub06_V_r_w = ( (|r_sys_processing_methodID) ? r_sub06_V_r_w : 1'h0 ) ;
	assign w_sub06_U_addr = ( (|r_sys_processing_methodID) ? r_sub06_U_addr : 9'sh0 ) ;
	assign w_sub06_U_datain = ( (|r_sys_processing_methodID) ? r_sub06_U_datain : 32'h0 ) ;
	assign w_sub06_U_r_w = ( (|r_sys_processing_methodID) ? r_sub06_U_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 9'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub05_T_addr = ( (|r_sys_processing_methodID) ? r_sub05_T_addr : 9'sh0 ) ;
	assign w_sub05_T_datain = ( (|r_sys_processing_methodID) ? r_sub05_T_datain : 32'h0 ) ;
	assign w_sub05_T_r_w = ( (|r_sys_processing_methodID) ? r_sub05_T_r_w : 1'h0 ) ;
	assign w_sub05_V_addr = ( (|r_sys_processing_methodID) ? r_sub05_V_addr : 9'sh0 ) ;
	assign w_sub05_V_datain = ( (|r_sys_processing_methodID) ? r_sub05_V_datain : 32'h0 ) ;
	assign w_sub05_V_r_w = ( (|r_sys_processing_methodID) ? r_sub05_V_r_w : 1'h0 ) ;
	assign w_sub05_U_addr = ( (|r_sys_processing_methodID) ? r_sub05_U_addr : 9'sh0 ) ;
	assign w_sub05_U_datain = ( (|r_sys_processing_methodID) ? r_sub05_U_datain : 32'h0 ) ;
	assign w_sub05_U_r_w = ( (|r_sys_processing_methodID) ? r_sub05_U_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 9'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_T_addr = ( (|r_sys_processing_methodID) ? r_sub04_T_addr : 9'sh0 ) ;
	assign w_sub04_T_datain = ( (|r_sys_processing_methodID) ? r_sub04_T_datain : 32'h0 ) ;
	assign w_sub04_T_r_w = ( (|r_sys_processing_methodID) ? r_sub04_T_r_w : 1'h0 ) ;
	assign w_sub04_V_addr = ( (|r_sys_processing_methodID) ? r_sub04_V_addr : 9'sh0 ) ;
	assign w_sub04_V_datain = ( (|r_sys_processing_methodID) ? r_sub04_V_datain : 32'h0 ) ;
	assign w_sub04_V_r_w = ( (|r_sys_processing_methodID) ? r_sub04_V_r_w : 1'h0 ) ;
	assign w_sub04_U_addr = ( (|r_sys_processing_methodID) ? r_sub04_U_addr : 9'sh0 ) ;
	assign w_sub04_U_datain = ( (|r_sys_processing_methodID) ? r_sub04_U_datain : 32'h0 ) ;
	assign w_sub04_U_r_w = ( (|r_sys_processing_methodID) ? r_sub04_U_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 9'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000080;
	assign w_sys_tmp3 = 32'sh00000081;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'h3d000000;
	assign w_sys_tmp7 = 32'h3c000000;
	assign w_sys_tmp8 = 32'h3c03126f;
	assign w_sys_tmp9 = 32'h3d03126f;
	assign w_sys_tmp10 = 32'h3f03126f;
	assign w_sys_tmp11 = 32'h4103126f;
	assign w_sys_tmp12 = ( !w_sys_tmp13 );
	assign w_sys_tmp13 = (r_run_my_16 < r_run_k_12);
	assign w_sys_tmp14 = (r_run_k_12 + w_sys_intOne);
	assign w_sys_tmp15 = ( !w_sys_tmp16 );
	assign w_sys_tmp16 = (r_run_mx_15 < r_run_j_13);
	assign w_sys_tmp18 = w_ip_MultFloat_product_0;
	assign w_sys_tmp19 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp20 = (r_run_k_12 - w_sys_intOne);
	assign w_sys_tmp22 = (w_sys_tmp23 + r_run_k_12);
	assign w_sys_tmp23 = (r_run_j_13 * w_sys_tmp24);
	assign w_sys_tmp24 = 32'sh00000081;
	assign w_sys_tmp25 = 32'h0;
	assign w_sys_tmp27 = (w_sys_tmp28 + r_run_k_12);
	assign w_sys_tmp28 = (r_run_copy2_j_30 * w_sys_tmp24);
	assign w_sys_tmp32 = (w_sys_tmp33 + r_run_k_12);
	assign w_sys_tmp33 = (r_run_copy1_j_29 * w_sys_tmp24);
	assign w_sys_tmp36 = 32'h42200000;
	assign w_sys_tmp37 = w_sys_tmp18;
	assign w_sys_tmp38 = 32'h3f800000;
	assign w_sys_tmp41 = (w_sys_tmp42 + r_run_k_12);
	assign w_sys_tmp42 = (r_run_copy0_j_28 * w_sys_tmp24);
	assign w_sys_tmp45 = (r_run_copy0_j_28 + w_sys_intOne);
	assign w_sys_tmp46 = (r_run_copy1_j_29 + w_sys_intOne);
	assign w_sys_tmp47 = (r_run_copy2_j_30 + w_sys_intOne);
	assign w_sys_tmp48 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp128 = r_sys_tmp4_float;
	assign w_sys_tmp226 = ( !w_sys_tmp227 );
	assign w_sys_tmp227 = (w_sys_tmp228 < r_run_k_12);
	assign w_sys_tmp228 = 32'sh00000041;
	assign w_sys_tmp229 = (r_run_k_12 + w_sys_intOne);
	assign w_sys_tmp230 = ( !w_sys_tmp231 );
	assign w_sys_tmp231 = (w_sys_tmp232 < r_run_j_13);
	assign w_sys_tmp232 = 32'sh00000021;
	assign w_sys_tmp235 = (w_sys_tmp236 + r_run_k_12);
	assign w_sys_tmp236 = (r_run_j_13 * w_sys_tmp237);
	assign w_sys_tmp237 = 32'sh00000081;
	assign w_sys_tmp238 = w_fld_U_2_dataout_1;
	assign w_sys_tmp239 = (w_sys_tmp240 + r_run_k_12);
	assign w_sys_tmp240 = (r_run_copy4_j_35 * w_sys_tmp237);
	assign w_sys_tmp243 = (w_sys_tmp244 + r_run_k_12);
	assign w_sys_tmp244 = (r_run_copy3_j_34 * w_sys_tmp237);
	assign w_sys_tmp246 = w_fld_V_3_dataout_1;
	assign w_sys_tmp247 = (w_sys_tmp248 + r_run_k_12);
	assign w_sys_tmp248 = (r_run_copy2_j_33 * w_sys_tmp237);
	assign w_sys_tmp251 = (w_sys_tmp252 + r_run_k_12);
	assign w_sys_tmp252 = (r_run_copy1_j_32 * w_sys_tmp237);
	assign w_sys_tmp254 = w_fld_T_0_dataout_1;
	assign w_sys_tmp255 = (w_sys_tmp256 + r_run_k_12);
	assign w_sys_tmp256 = (r_run_copy0_j_31 * w_sys_tmp237);
	assign w_sys_tmp258 = (r_run_copy0_j_31 + w_sys_intOne);
	assign w_sys_tmp259 = (r_run_copy1_j_32 + w_sys_intOne);
	assign w_sys_tmp260 = (r_run_copy2_j_33 + w_sys_intOne);
	assign w_sys_tmp261 = (r_run_copy3_j_34 + w_sys_intOne);
	assign w_sys_tmp262 = (r_run_copy4_j_35 + w_sys_intOne);
	assign w_sys_tmp263 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp444 = 32'sh00000020;
	assign w_sys_tmp445 = ( !w_sys_tmp446 );
	assign w_sys_tmp446 = (w_sys_tmp447 < r_run_j_13);
	assign w_sys_tmp447 = 32'sh00000041;
	assign w_sys_tmp450 = (w_sys_tmp451 + r_run_k_12);
	assign w_sys_tmp451 = (r_run_j_13 * w_sys_tmp452);
	assign w_sys_tmp452 = 32'sh00000081;
	assign w_sys_tmp453 = w_fld_U_2_dataout_1;
	assign w_sys_tmp454 = (w_sys_tmp455 + r_run_k_12);
	assign w_sys_tmp455 = (r_run_copy4_j_40 * w_sys_tmp452);
	assign w_sys_tmp458 = (w_sys_tmp459 + r_run_k_12);
	assign w_sys_tmp459 = (r_run_copy3_j_39 * w_sys_tmp452);
	assign w_sys_tmp461 = w_fld_V_3_dataout_1;
	assign w_sys_tmp462 = (w_sys_tmp463 + r_run_k_12);
	assign w_sys_tmp463 = (r_run_copy2_j_38 * w_sys_tmp452);
	assign w_sys_tmp466 = (w_sys_tmp467 + r_run_k_12);
	assign w_sys_tmp467 = (r_run_copy1_j_37 * w_sys_tmp452);
	assign w_sys_tmp469 = w_fld_T_0_dataout_1;
	assign w_sys_tmp470 = (w_sys_tmp471 + r_run_k_12);
	assign w_sys_tmp471 = (r_run_copy0_j_36 * w_sys_tmp452);
	assign w_sys_tmp473 = (r_run_copy0_j_36 + w_sys_intOne);
	assign w_sys_tmp474 = (r_run_copy1_j_37 + w_sys_intOne);
	assign w_sys_tmp475 = (r_run_copy2_j_38 + w_sys_intOne);
	assign w_sys_tmp476 = (r_run_copy3_j_39 + w_sys_intOne);
	assign w_sys_tmp477 = (r_run_copy4_j_40 + w_sys_intOne);
	assign w_sys_tmp478 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp659 = 32'sh00000040;
	assign w_sys_tmp660 = ( !w_sys_tmp661 );
	assign w_sys_tmp661 = (w_sys_tmp662 < r_run_j_13);
	assign w_sys_tmp662 = 32'sh00000061;
	assign w_sys_tmp665 = (w_sys_tmp666 + r_run_k_12);
	assign w_sys_tmp666 = (r_run_j_13 * w_sys_tmp667);
	assign w_sys_tmp667 = 32'sh00000081;
	assign w_sys_tmp668 = w_fld_U_2_dataout_1;
	assign w_sys_tmp669 = (w_sys_tmp670 + r_run_k_12);
	assign w_sys_tmp670 = (r_run_copy4_j_45 * w_sys_tmp667);
	assign w_sys_tmp673 = (w_sys_tmp674 + r_run_k_12);
	assign w_sys_tmp674 = (r_run_copy3_j_44 * w_sys_tmp667);
	assign w_sys_tmp676 = w_fld_V_3_dataout_1;
	assign w_sys_tmp677 = (w_sys_tmp678 + r_run_k_12);
	assign w_sys_tmp678 = (r_run_copy2_j_43 * w_sys_tmp667);
	assign w_sys_tmp681 = (w_sys_tmp682 + r_run_k_12);
	assign w_sys_tmp682 = (r_run_copy1_j_42 * w_sys_tmp667);
	assign w_sys_tmp684 = w_fld_T_0_dataout_1;
	assign w_sys_tmp685 = (w_sys_tmp686 + r_run_k_12);
	assign w_sys_tmp686 = (r_run_copy0_j_41 * w_sys_tmp667);
	assign w_sys_tmp688 = (r_run_copy0_j_41 + w_sys_intOne);
	assign w_sys_tmp689 = (r_run_copy1_j_42 + w_sys_intOne);
	assign w_sys_tmp690 = (r_run_copy2_j_43 + w_sys_intOne);
	assign w_sys_tmp691 = (r_run_copy3_j_44 + w_sys_intOne);
	assign w_sys_tmp692 = (r_run_copy4_j_45 + w_sys_intOne);
	assign w_sys_tmp693 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp874 = 32'sh00000060;
	assign w_sys_tmp875 = ( !w_sys_tmp876 );
	assign w_sys_tmp876 = (w_sys_tmp877 < r_run_j_13);
	assign w_sys_tmp877 = 32'sh00000081;
	assign w_sys_tmp880 = (w_sys_tmp881 + r_run_k_12);
	assign w_sys_tmp881 = (r_run_j_13 * w_sys_tmp882);
	assign w_sys_tmp882 = 32'sh00000081;
	assign w_sys_tmp883 = w_fld_U_2_dataout_1;
	assign w_sys_tmp884 = (w_sys_tmp885 + r_run_k_12);
	assign w_sys_tmp885 = (r_run_copy4_j_50 * w_sys_tmp882);
	assign w_sys_tmp888 = (w_sys_tmp889 + r_run_k_12);
	assign w_sys_tmp889 = (r_run_copy3_j_49 * w_sys_tmp882);
	assign w_sys_tmp891 = w_fld_V_3_dataout_1;
	assign w_sys_tmp892 = (w_sys_tmp893 + r_run_k_12);
	assign w_sys_tmp893 = (r_run_copy2_j_48 * w_sys_tmp882);
	assign w_sys_tmp896 = (w_sys_tmp897 + r_run_k_12);
	assign w_sys_tmp897 = (r_run_copy1_j_47 * w_sys_tmp882);
	assign w_sys_tmp899 = w_fld_T_0_dataout_1;
	assign w_sys_tmp900 = (w_sys_tmp901 + r_run_k_12);
	assign w_sys_tmp901 = (r_run_copy0_j_46 * w_sys_tmp882);
	assign w_sys_tmp903 = (r_run_copy0_j_46 + w_sys_intOne);
	assign w_sys_tmp904 = (r_run_copy1_j_47 + w_sys_intOne);
	assign w_sys_tmp905 = (r_run_copy2_j_48 + w_sys_intOne);
	assign w_sys_tmp906 = (r_run_copy3_j_49 + w_sys_intOne);
	assign w_sys_tmp907 = (r_run_copy4_j_50 + w_sys_intOne);
	assign w_sys_tmp908 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp1089 = 32'sh00000040;
	assign w_sys_tmp1090 = ( !w_sys_tmp1091 );
	assign w_sys_tmp1091 = (w_sys_tmp1092 < r_run_k_12);
	assign w_sys_tmp1092 = 32'sh00000081;
	assign w_sys_tmp1093 = (r_run_k_12 + w_sys_intOne);
	assign w_sys_tmp1094 = ( !w_sys_tmp1095 );
	assign w_sys_tmp1095 = (w_sys_tmp1096 < r_run_j_13);
	assign w_sys_tmp1096 = 32'sh00000021;
	assign w_sys_tmp1099 = (w_sys_tmp1100 + r_run_k_12);
	assign w_sys_tmp1100 = (r_run_j_13 * w_sys_tmp1101);
	assign w_sys_tmp1101 = 32'sh00000081;
	assign w_sys_tmp1102 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1103 = (w_sys_tmp1104 + r_run_k_12);
	assign w_sys_tmp1104 = (r_run_copy4_j_55 * w_sys_tmp1101);
	assign w_sys_tmp1107 = (w_sys_tmp1108 + r_run_k_12);
	assign w_sys_tmp1108 = (r_run_copy3_j_54 * w_sys_tmp1101);
	assign w_sys_tmp1110 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1111 = (w_sys_tmp1112 + r_run_k_12);
	assign w_sys_tmp1112 = (r_run_copy2_j_53 * w_sys_tmp1101);
	assign w_sys_tmp1115 = (w_sys_tmp1116 + r_run_k_12);
	assign w_sys_tmp1116 = (r_run_copy1_j_52 * w_sys_tmp1101);
	assign w_sys_tmp1118 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1119 = (w_sys_tmp1120 + r_run_k_12);
	assign w_sys_tmp1120 = (r_run_copy0_j_51 * w_sys_tmp1101);
	assign w_sys_tmp1122 = (r_run_copy0_j_51 + w_sys_intOne);
	assign w_sys_tmp1123 = (r_run_copy1_j_52 + w_sys_intOne);
	assign w_sys_tmp1124 = (r_run_copy2_j_53 + w_sys_intOne);
	assign w_sys_tmp1125 = (r_run_copy3_j_54 + w_sys_intOne);
	assign w_sys_tmp1126 = (r_run_copy4_j_55 + w_sys_intOne);
	assign w_sys_tmp1127 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp1308 = 32'sh00000020;
	assign w_sys_tmp1309 = ( !w_sys_tmp1310 );
	assign w_sys_tmp1310 = (w_sys_tmp1311 < r_run_j_13);
	assign w_sys_tmp1311 = 32'sh00000041;
	assign w_sys_tmp1314 = (w_sys_tmp1315 + r_run_k_12);
	assign w_sys_tmp1315 = (r_run_j_13 * w_sys_tmp1316);
	assign w_sys_tmp1316 = 32'sh00000081;
	assign w_sys_tmp1317 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1318 = (w_sys_tmp1319 + r_run_k_12);
	assign w_sys_tmp1319 = (r_run_copy4_j_60 * w_sys_tmp1316);
	assign w_sys_tmp1322 = (w_sys_tmp1323 + r_run_k_12);
	assign w_sys_tmp1323 = (r_run_copy3_j_59 * w_sys_tmp1316);
	assign w_sys_tmp1325 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1326 = (w_sys_tmp1327 + r_run_k_12);
	assign w_sys_tmp1327 = (r_run_copy2_j_58 * w_sys_tmp1316);
	assign w_sys_tmp1330 = (w_sys_tmp1331 + r_run_k_12);
	assign w_sys_tmp1331 = (r_run_copy1_j_57 * w_sys_tmp1316);
	assign w_sys_tmp1333 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1334 = (w_sys_tmp1335 + r_run_k_12);
	assign w_sys_tmp1335 = (r_run_copy0_j_56 * w_sys_tmp1316);
	assign w_sys_tmp1337 = (r_run_copy0_j_56 + w_sys_intOne);
	assign w_sys_tmp1338 = (r_run_copy1_j_57 + w_sys_intOne);
	assign w_sys_tmp1339 = (r_run_copy2_j_58 + w_sys_intOne);
	assign w_sys_tmp1340 = (r_run_copy3_j_59 + w_sys_intOne);
	assign w_sys_tmp1341 = (r_run_copy4_j_60 + w_sys_intOne);
	assign w_sys_tmp1342 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp1523 = 32'sh00000040;
	assign w_sys_tmp1524 = ( !w_sys_tmp1525 );
	assign w_sys_tmp1525 = (w_sys_tmp1526 < r_run_j_13);
	assign w_sys_tmp1526 = 32'sh00000061;
	assign w_sys_tmp1529 = (w_sys_tmp1530 + r_run_k_12);
	assign w_sys_tmp1530 = (r_run_j_13 * w_sys_tmp1531);
	assign w_sys_tmp1531 = 32'sh00000081;
	assign w_sys_tmp1532 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1533 = (w_sys_tmp1534 + r_run_k_12);
	assign w_sys_tmp1534 = (r_run_copy4_j_65 * w_sys_tmp1531);
	assign w_sys_tmp1537 = (w_sys_tmp1538 + r_run_k_12);
	assign w_sys_tmp1538 = (r_run_copy3_j_64 * w_sys_tmp1531);
	assign w_sys_tmp1540 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1541 = (w_sys_tmp1542 + r_run_k_12);
	assign w_sys_tmp1542 = (r_run_copy2_j_63 * w_sys_tmp1531);
	assign w_sys_tmp1545 = (w_sys_tmp1546 + r_run_k_12);
	assign w_sys_tmp1546 = (r_run_copy1_j_62 * w_sys_tmp1531);
	assign w_sys_tmp1548 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1549 = (w_sys_tmp1550 + r_run_k_12);
	assign w_sys_tmp1550 = (r_run_copy0_j_61 * w_sys_tmp1531);
	assign w_sys_tmp1552 = (r_run_copy0_j_61 + w_sys_intOne);
	assign w_sys_tmp1553 = (r_run_copy1_j_62 + w_sys_intOne);
	assign w_sys_tmp1554 = (r_run_copy2_j_63 + w_sys_intOne);
	assign w_sys_tmp1555 = (r_run_copy3_j_64 + w_sys_intOne);
	assign w_sys_tmp1556 = (r_run_copy4_j_65 + w_sys_intOne);
	assign w_sys_tmp1557 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp1738 = 32'sh00000060;
	assign w_sys_tmp1739 = ( !w_sys_tmp1740 );
	assign w_sys_tmp1740 = (w_sys_tmp1741 < r_run_j_13);
	assign w_sys_tmp1741 = 32'sh00000081;
	assign w_sys_tmp1744 = (w_sys_tmp1745 + r_run_k_12);
	assign w_sys_tmp1745 = (r_run_j_13 * w_sys_tmp1746);
	assign w_sys_tmp1746 = 32'sh00000081;
	assign w_sys_tmp1747 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1748 = (w_sys_tmp1749 + r_run_k_12);
	assign w_sys_tmp1749 = (r_run_copy4_j_70 * w_sys_tmp1746);
	assign w_sys_tmp1752 = (w_sys_tmp1753 + r_run_k_12);
	assign w_sys_tmp1753 = (r_run_copy3_j_69 * w_sys_tmp1746);
	assign w_sys_tmp1755 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1756 = (w_sys_tmp1757 + r_run_k_12);
	assign w_sys_tmp1757 = (r_run_copy2_j_68 * w_sys_tmp1746);
	assign w_sys_tmp1760 = (w_sys_tmp1761 + r_run_k_12);
	assign w_sys_tmp1761 = (r_run_copy1_j_67 * w_sys_tmp1746);
	assign w_sys_tmp1763 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1764 = (w_sys_tmp1765 + r_run_k_12);
	assign w_sys_tmp1765 = (r_run_copy0_j_66 * w_sys_tmp1746);
	assign w_sys_tmp1767 = (r_run_copy0_j_66 + w_sys_intOne);
	assign w_sys_tmp1768 = (r_run_copy1_j_67 + w_sys_intOne);
	assign w_sys_tmp1769 = (r_run_copy2_j_68 + w_sys_intOne);
	assign w_sys_tmp1770 = (r_run_copy3_j_69 + w_sys_intOne);
	assign w_sys_tmp1771 = (r_run_copy4_j_70 + w_sys_intOne);
	assign w_sys_tmp1772 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp1953 = ( !w_sys_tmp1954 );
	assign w_sys_tmp1954 = (r_run_nlast_27 < r_run_n_14);
	assign w_sys_tmp1955 = (r_run_n_14 + w_sys_intOne);
	assign w_sys_tmp1956 = 32'sh00000002;
	assign w_sys_tmp1957 = ( !w_sys_tmp1958 );
	assign w_sys_tmp1958 = (w_sys_tmp1959 < r_run_k_12);
	assign w_sys_tmp1959 = 32'sh00000040;
	assign w_sys_tmp1962 = (w_sys_tmp1963 + r_run_k_12);
	assign w_sys_tmp1963 = 32'sh000010a1;
	assign w_sys_tmp1964 = w_sub01_result_dataout;
	assign w_sys_tmp1968 = (w_sys_tmp1969 + r_run_k_12);
	assign w_sys_tmp1969 = 32'sh00003060;
	assign w_sys_tmp1970 = w_sub02_result_dataout;
	assign w_sys_tmp1974 = (w_sys_tmp1975 + r_run_k_12);
	assign w_sys_tmp1975 = 32'sh00002040;
	assign w_sys_tmp1976 = w_sub00_result_dataout;
	assign w_sys_tmp1980 = (w_sys_tmp1981 + r_run_k_12);
	assign w_sys_tmp1981 = 32'sh000030e1;
	assign w_sys_tmp1985 = (w_sys_tmp1986 + r_run_k_12);
	assign w_sys_tmp1986 = 32'sh00001020;
	assign w_sys_tmp1990 = (w_sys_tmp1991 + r_run_k_12);
	assign w_sys_tmp1991 = 32'sh000020c1;
	assign w_sys_tmp1994 = (r_run_k_12 + w_sys_intOne);
	assign w_sys_tmp1995 = 32'sh00000002;
	assign w_sys_tmp1996 = ( !w_sys_tmp1997 );
	assign w_sys_tmp1997 = (w_sys_tmp1998 < r_run_j_13);
	assign w_sys_tmp1998 = 32'sh00000020;
	assign w_sys_tmp2001 = (w_sys_tmp2002 + w_sys_tmp2004);
	assign w_sys_tmp2002 = (r_run_j_13 * w_sys_tmp2003);
	assign w_sys_tmp2003 = 32'sh00000081;
	assign w_sys_tmp2004 = 32'sh00000041;
	assign w_sys_tmp2005 = w_sub04_result_dataout;
	assign w_sys_tmp2006 = (w_sys_tmp2007 + w_sys_tmp2004);
	assign w_sys_tmp2007 = (r_run_copy2_j_73 * w_sys_tmp2003);
	assign w_sys_tmp2011 = (w_sys_tmp2012 + w_sys_tmp2014);
	assign w_sys_tmp2012 = (r_run_copy1_j_72 * w_sys_tmp2003);
	assign w_sys_tmp2014 = 32'sh00000040;
	assign w_sys_tmp2015 = w_sub00_result_dataout;
	assign w_sys_tmp2016 = (w_sys_tmp2017 + w_sys_tmp2014);
	assign w_sys_tmp2017 = (r_run_copy0_j_71 * w_sys_tmp2003);
	assign w_sys_tmp2020 = (r_run_copy0_j_71 + w_sys_intOne);
	assign w_sys_tmp2021 = (r_run_copy1_j_72 + w_sys_intOne);
	assign w_sys_tmp2022 = (r_run_copy2_j_73 + w_sys_intOne);
	assign w_sys_tmp2023 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp2168 = 32'sh00000021;
	assign w_sys_tmp2169 = ( !w_sys_tmp2170 );
	assign w_sys_tmp2170 = (w_sys_tmp2171 < r_run_j_13);
	assign w_sys_tmp2171 = 32'sh00000040;
	assign w_sys_tmp2174 = (w_sys_tmp2175 + w_sys_tmp2177);
	assign w_sys_tmp2175 = (r_run_j_13 * w_sys_tmp2176);
	assign w_sys_tmp2176 = 32'sh00000081;
	assign w_sys_tmp2177 = 32'sh00000041;
	assign w_sys_tmp2178 = w_sub05_result_dataout;
	assign w_sys_tmp2179 = (w_sys_tmp2180 + w_sys_tmp2177);
	assign w_sys_tmp2180 = (r_run_copy2_j_76 * w_sys_tmp2176);
	assign w_sys_tmp2184 = (w_sys_tmp2185 + w_sys_tmp2187);
	assign w_sys_tmp2185 = (r_run_copy1_j_75 * w_sys_tmp2176);
	assign w_sys_tmp2187 = 32'sh00000040;
	assign w_sys_tmp2188 = w_sub01_result_dataout;
	assign w_sys_tmp2189 = (w_sys_tmp2190 + w_sys_tmp2187);
	assign w_sys_tmp2190 = (r_run_copy0_j_74 * w_sys_tmp2176);
	assign w_sys_tmp2193 = (r_run_copy0_j_74 + w_sys_intOne);
	assign w_sys_tmp2194 = (r_run_copy1_j_75 + w_sys_intOne);
	assign w_sys_tmp2195 = (r_run_copy2_j_76 + w_sys_intOne);
	assign w_sys_tmp2196 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp2341 = 32'sh00000041;
	assign w_sys_tmp2342 = ( !w_sys_tmp2343 );
	assign w_sys_tmp2343 = (w_sys_tmp2344 < r_run_j_13);
	assign w_sys_tmp2344 = 32'sh00000060;
	assign w_sys_tmp2347 = (w_sys_tmp2348 + w_sys_tmp2350);
	assign w_sys_tmp2348 = (r_run_j_13 * w_sys_tmp2349);
	assign w_sys_tmp2349 = 32'sh00000081;
	assign w_sys_tmp2350 = 32'sh00000041;
	assign w_sys_tmp2351 = w_sub06_result_dataout;
	assign w_sys_tmp2352 = (w_sys_tmp2353 + w_sys_tmp2350);
	assign w_sys_tmp2353 = (r_run_copy2_j_79 * w_sys_tmp2349);
	assign w_sys_tmp2357 = (w_sys_tmp2358 + w_sys_tmp2360);
	assign w_sys_tmp2358 = (r_run_copy1_j_78 * w_sys_tmp2349);
	assign w_sys_tmp2360 = 32'sh00000040;
	assign w_sys_tmp2361 = w_sub02_result_dataout;
	assign w_sys_tmp2362 = (w_sys_tmp2363 + w_sys_tmp2360);
	assign w_sys_tmp2363 = (r_run_copy0_j_77 * w_sys_tmp2349);
	assign w_sys_tmp2366 = (r_run_copy0_j_77 + w_sys_intOne);
	assign w_sys_tmp2367 = (r_run_copy1_j_78 + w_sys_intOne);
	assign w_sys_tmp2368 = (r_run_copy2_j_79 + w_sys_intOne);
	assign w_sys_tmp2369 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp2514 = 32'sh00000061;
	assign w_sys_tmp2515 = ( !w_sys_tmp2516 );
	assign w_sys_tmp2516 = (w_sys_tmp2517 < r_run_j_13);
	assign w_sys_tmp2517 = 32'sh00000080;
	assign w_sys_tmp2520 = (w_sys_tmp2521 + w_sys_tmp2523);
	assign w_sys_tmp2521 = (r_run_j_13 * w_sys_tmp2522);
	assign w_sys_tmp2522 = 32'sh00000081;
	assign w_sys_tmp2523 = 32'sh00000041;
	assign w_sys_tmp2524 = w_sub07_result_dataout;
	assign w_sys_tmp2525 = (w_sys_tmp2526 + w_sys_tmp2523);
	assign w_sys_tmp2526 = (r_run_copy2_j_82 * w_sys_tmp2522);
	assign w_sys_tmp2530 = (w_sys_tmp2531 + w_sys_tmp2533);
	assign w_sys_tmp2531 = (r_run_copy1_j_81 * w_sys_tmp2522);
	assign w_sys_tmp2533 = 32'sh00000040;
	assign w_sys_tmp2534 = w_sub03_result_dataout;
	assign w_sys_tmp2535 = (w_sys_tmp2536 + w_sys_tmp2533);
	assign w_sys_tmp2536 = (r_run_copy0_j_80 * w_sys_tmp2522);
	assign w_sys_tmp2539 = (r_run_copy0_j_80 + w_sys_intOne);
	assign w_sys_tmp2540 = (r_run_copy1_j_81 + w_sys_intOne);
	assign w_sys_tmp2541 = (r_run_copy2_j_82 + w_sys_intOne);
	assign w_sys_tmp2542 = (r_run_j_13 + w_sys_intOne);
	assign w_sys_tmp2687 = 32'sh00000041;
	assign w_sys_tmp2688 = ( !w_sys_tmp2689 );
	assign w_sys_tmp2689 = (w_sys_tmp2690 < r_run_k_12);
	assign w_sys_tmp2690 = 32'sh00000080;
	assign w_sys_tmp2693 = (w_sys_tmp2694 + r_run_k_12);
	assign w_sys_tmp2694 = 32'sh000010a1;
	assign w_sys_tmp2695 = w_sub05_result_dataout;
	assign w_sys_tmp2699 = (w_sys_tmp2700 + r_run_k_12);
	assign w_sys_tmp2700 = 32'sh00001020;
	assign w_sys_tmp2701 = w_sub04_result_dataout;
	assign w_sys_tmp2705 = (w_sys_tmp2706 + r_run_k_12);
	assign w_sys_tmp2706 = 32'sh000020c1;
	assign w_sys_tmp2710 = (w_sys_tmp2711 + r_run_k_12);
	assign w_sys_tmp2711 = 32'sh00003060;
	assign w_sys_tmp2712 = w_sub06_result_dataout;
	assign w_sys_tmp2716 = (w_sys_tmp2717 + r_run_k_12);
	assign w_sys_tmp2717 = 32'sh00002040;
	assign w_sys_tmp2722 = (w_sys_tmp2723 + r_run_k_12);
	assign w_sys_tmp2723 = 32'sh000030e1;
	assign w_sys_tmp2726 = (r_run_k_12 + w_sys_intOne);


	sub03
		sub03_inst(
			.i_fld_T_0_addr_0 (w_sub03_T_addr),
			.i_fld_T_0_datain_0 (w_sub03_T_datain),
			.o_fld_T_0_dataout_0 (w_sub03_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub03_T_r_w),
			.i_fld_U_2_addr_0 (w_sub03_U_addr),
			.i_fld_U_2_datain_0 (w_sub03_U_datain),
			.o_fld_U_2_dataout_0 (w_sub03_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub03_U_r_w),
			.i_fld_V_1_addr_0 (w_sub03_V_addr),
			.i_fld_V_1_datain_0 (w_sub03_V_datain),
			.o_fld_V_1_dataout_0 (w_sub03_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub03_V_r_w),
			.i_fld_result_3_addr_0 (w_sub03_result_addr),
			.i_fld_result_3_datain_0 (w_sub03_result_datain),
			.o_fld_result_3_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub03_result_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_T_0_addr_0 (w_sub02_T_addr),
			.i_fld_T_0_datain_0 (w_sub02_T_datain),
			.o_fld_T_0_dataout_0 (w_sub02_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub02_T_r_w),
			.i_fld_U_2_addr_0 (w_sub02_U_addr),
			.i_fld_U_2_datain_0 (w_sub02_U_datain),
			.o_fld_U_2_dataout_0 (w_sub02_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub02_U_r_w),
			.i_fld_V_1_addr_0 (w_sub02_V_addr),
			.i_fld_V_1_datain_0 (w_sub02_V_datain),
			.o_fld_V_1_dataout_0 (w_sub02_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub02_V_r_w),
			.i_fld_result_3_addr_0 (w_sub02_result_addr),
			.i_fld_result_3_datain_0 (w_sub02_result_datain),
			.o_fld_result_3_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub02_result_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_T_0_addr_0 (w_sub01_T_addr),
			.i_fld_T_0_datain_0 (w_sub01_T_datain),
			.o_fld_T_0_dataout_0 (w_sub01_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub01_T_r_w),
			.i_fld_U_2_addr_0 (w_sub01_U_addr),
			.i_fld_U_2_datain_0 (w_sub01_U_datain),
			.o_fld_U_2_dataout_0 (w_sub01_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub01_U_r_w),
			.i_fld_V_1_addr_0 (w_sub01_V_addr),
			.i_fld_V_1_datain_0 (w_sub01_V_datain),
			.o_fld_V_1_dataout_0 (w_sub01_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub01_V_r_w),
			.i_fld_result_3_addr_0 (w_sub01_result_addr),
			.i_fld_result_3_datain_0 (w_sub01_result_datain),
			.o_fld_result_3_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub01_result_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_T_0_addr_0 (w_sub00_T_addr),
			.i_fld_T_0_datain_0 (w_sub00_T_datain),
			.o_fld_T_0_dataout_0 (w_sub00_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub00_T_r_w),
			.i_fld_U_2_addr_0 (w_sub00_U_addr),
			.i_fld_U_2_datain_0 (w_sub00_U_datain),
			.o_fld_U_2_dataout_0 (w_sub00_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub00_U_r_w),
			.i_fld_V_1_addr_0 (w_sub00_V_addr),
			.i_fld_V_1_datain_0 (w_sub00_V_datain),
			.o_fld_V_1_dataout_0 (w_sub00_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub00_V_r_w),
			.i_fld_result_3_addr_0 (w_sub00_result_addr),
			.i_fld_result_3_datain_0 (w_sub00_result_datain),
			.o_fld_result_3_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub00_result_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_T_0_addr_0 (w_sub07_T_addr),
			.i_fld_T_0_datain_0 (w_sub07_T_datain),
			.o_fld_T_0_dataout_0 (w_sub07_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub07_T_r_w),
			.i_fld_U_2_addr_0 (w_sub07_U_addr),
			.i_fld_U_2_datain_0 (w_sub07_U_datain),
			.o_fld_U_2_dataout_0 (w_sub07_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub07_U_r_w),
			.i_fld_V_1_addr_0 (w_sub07_V_addr),
			.i_fld_V_1_datain_0 (w_sub07_V_datain),
			.o_fld_V_1_dataout_0 (w_sub07_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub07_V_r_w),
			.i_fld_result_3_addr_0 (w_sub07_result_addr),
			.i_fld_result_3_datain_0 (w_sub07_result_datain),
			.o_fld_result_3_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub07_result_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_T_0_addr_0 (w_sub06_T_addr),
			.i_fld_T_0_datain_0 (w_sub06_T_datain),
			.o_fld_T_0_dataout_0 (w_sub06_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub06_T_r_w),
			.i_fld_U_2_addr_0 (w_sub06_U_addr),
			.i_fld_U_2_datain_0 (w_sub06_U_datain),
			.o_fld_U_2_dataout_0 (w_sub06_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub06_U_r_w),
			.i_fld_V_1_addr_0 (w_sub06_V_addr),
			.i_fld_V_1_datain_0 (w_sub06_V_datain),
			.o_fld_V_1_dataout_0 (w_sub06_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub06_V_r_w),
			.i_fld_result_3_addr_0 (w_sub06_result_addr),
			.i_fld_result_3_datain_0 (w_sub06_result_datain),
			.o_fld_result_3_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub06_result_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_T_0_addr_0 (w_sub05_T_addr),
			.i_fld_T_0_datain_0 (w_sub05_T_datain),
			.o_fld_T_0_dataout_0 (w_sub05_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub05_T_r_w),
			.i_fld_U_2_addr_0 (w_sub05_U_addr),
			.i_fld_U_2_datain_0 (w_sub05_U_datain),
			.o_fld_U_2_dataout_0 (w_sub05_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub05_U_r_w),
			.i_fld_V_1_addr_0 (w_sub05_V_addr),
			.i_fld_V_1_datain_0 (w_sub05_V_datain),
			.o_fld_V_1_dataout_0 (w_sub05_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub05_V_r_w),
			.i_fld_result_3_addr_0 (w_sub05_result_addr),
			.i_fld_result_3_datain_0 (w_sub05_result_datain),
			.o_fld_result_3_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub05_result_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_T_0_addr_0 (w_sub04_T_addr),
			.i_fld_T_0_datain_0 (w_sub04_T_datain),
			.o_fld_T_0_dataout_0 (w_sub04_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub04_T_r_w),
			.i_fld_U_2_addr_0 (w_sub04_U_addr),
			.i_fld_U_2_datain_0 (w_sub04_U_datain),
			.o_fld_U_2_dataout_0 (w_sub04_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub04_U_r_w),
			.i_fld_V_1_addr_0 (w_sub04_V_addr),
			.i_fld_V_1_datain_0 (w_sub04_V_datain),
			.o_fld_V_1_dataout_0 (w_sub04_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub04_V_r_w),
			.i_fld_result_3_addr_0 (w_sub04_result_addr),
			.i_fld_result_3_datain_0 (w_sub04_result_datain),
			.o_fld_result_3_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub04_result_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_V_3(
			.clk (clock),
			.ce_0 (w_fld_V_3_ce_0),
			.addr_0 (w_fld_V_3_addr_0),
			.datain_0 (w_fld_V_3_datain_0),
			.dataout_0 (w_fld_V_3_dataout_0),
			.r_w_0 (w_fld_V_3_r_w_0),
			.ce_1 (w_fld_V_3_ce_1),
			.addr_1 (r_fld_V_3_addr_1),
			.datain_1 (r_fld_V_3_datain_1),
			.dataout_1 (w_fld_V_3_dataout_1),
			.r_w_1 (r_fld_V_3_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp38;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h7<=r_sys_run_step && r_sys_run_step<=6'hb) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'hf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_19;

									end
									else
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h16)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp36;

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp18;

									end
									else
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h18)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h7<=r_sys_run_step && r_sys_run_step<=6'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp37;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h16)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h75: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp15) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp226) ? 7'h14 : 7'h2c);

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h15;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp230) ? 7'h18 : 7'h1a);

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 7'h15;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp445) ? 7'h1e : 7'h20);

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp660) ? 7'h24 : 7'h26);

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp875) ? 7'h2a : 7'h11);

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1090) ? 7'h31 : 7'h49);

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h32;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1094) ? 7'h35 : 7'h37);

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 7'h32;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h38;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1309) ? 7'h3b : 7'h3d);

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 7'h38;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h3e;

									end
								end

							endcase
						end

						7'h3e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1524) ? 7'h41 : 7'h43);

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 7'h3e;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h44;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1739) ? 7'h47 : 7'h2e);

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 7'h44;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h4a;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1953) ? 7'h4d : 7'h75);

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h4a;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 7'h4f;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_run_stage) 
								4'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 7'h51;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h52;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1957) ? 7'h55 : 7'h57);

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 7'h52;

									end
								end

							endcase
						end

						7'h57: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h58;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1996) ? 7'h5b : 7'h5d);

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_phase <= 7'h58;

									end
								end

							endcase
						end

						7'h5d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h5e;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2169) ? 7'h61 : 7'h63);

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_phase <= 7'h5e;

									end
								end

							endcase
						end

						7'h63: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h64;

									end
								end

							endcase
						end

						7'h64: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2342) ? 7'h67 : 7'h69);

									end
								end

							endcase
						end

						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_phase <= 7'h64;

									end
								end

							endcase
						end

						7'h69: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h6a;

									end
								end

							endcase
						end

						7'h6a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2515) ? 7'h6d : 7'h6f);

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_phase <= 7'h6a;

									end
								end

							endcase
						end

						7'h6f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 7'h70;

									end
								end

							endcase
						end

						7'h70: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2688) ? 7'h73 : 7'h4b);

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sys_run_phase <= 7'h70;

									end
								end

							endcase
						end

						7'h75: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h3e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h57: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h5d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h63: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h64: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h69: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h6a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h6f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h70: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h3e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h57: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h28)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h5d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h28)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h63: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h64: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h28)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h69: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h6a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h28)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h29)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h6f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h70: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h9)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h75: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp22[14:0] );

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp255[14:0] );

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp470[14:0] );

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp685[14:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp900[14:0] );

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1119[14:0] );

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1334[14:0] );

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1549[14:0] );

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1764[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp27[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h75: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp32[14:0] );

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp239[14:0] );

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp454[14:0] );

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp669[14:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp884[14:0] );

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1103[14:0] );

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1318[14:0] );

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1533[14:0] );

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1748[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp41[14:0] );

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp247[14:0] );

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp462[14:0] );

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp677[14:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp892[14:0] );

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1111[14:0] );

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1326[14:0] );

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1541[14:0] );

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1756[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_fld_V_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_12 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_12 <= w_sys_tmp14;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_12 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_12 <= w_sys_tmp229;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_12 <= w_sys_tmp1089;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_12 <= w_sys_tmp1093;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_12 <= w_sys_tmp1956;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_run_k_12 <= w_sys_tmp1994;

									end
								end

							endcase
						end

						7'h6f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_12 <= w_sys_tmp2687;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_run_k_12 <= w_sys_tmp2726;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_13 <= w_sys_tmp48;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_13 <= w_sys_tmp263;

									end
								end

							endcase
						end

						7'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_tmp444;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_13 <= w_sys_tmp478;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_tmp659;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_13 <= w_sys_tmp693;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_tmp874;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_13 <= w_sys_tmp908;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_13 <= w_sys_tmp1127;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_tmp1308;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_13 <= w_sys_tmp1342;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_tmp1523;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_13 <= w_sys_tmp1557;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_tmp1738;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_13 <= w_sys_tmp1772;

									end
								end

							endcase
						end

						7'h57: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_tmp1995;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_run_j_13 <= w_sys_tmp2023;

									end
								end

							endcase
						end

						7'h5d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_tmp2168;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_run_j_13 <= w_sys_tmp2196;

									end
								end

							endcase
						end

						7'h63: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_tmp2341;

									end
								end

							endcase
						end

						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_run_j_13 <= w_sys_tmp2369;

									end
								end

							endcase
						end

						7'h69: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_13 <= w_sys_tmp2514;

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_run_j_13 <= w_sys_tmp2542;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h49: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_14 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_14 <= w_sys_tmp1955;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_mx_15 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_my_16 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dt_17 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dx_18 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dy_19 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r1_20 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r2_21 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r3_22 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r4_23 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14)) begin
										r_run_YY_24 <= w_sys_tmp18;

									end
									else
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h11)) begin
										r_run_YY_24 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_kx_25 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_ky_26 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_nlast_27 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_28 <= r_run_j_13;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_28 <= w_sys_tmp45;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_29 <= r_run_j_13;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_run_copy1_j_29 <= w_sys_tmp46;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_30 <= r_run_j_13;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_30 <= w_sys_tmp47;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_31 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_31 <= w_sys_tmp258;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_32 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_32 <= w_sys_tmp259;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_33 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_33 <= w_sys_tmp260;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_34 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_34 <= w_sys_tmp261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_35 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_35 <= w_sys_tmp262;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1a: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_36 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_36 <= w_sys_tmp473;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1a: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_37 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_37 <= w_sys_tmp474;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1a: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_38 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_38 <= w_sys_tmp475;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1a: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_39 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_39 <= w_sys_tmp476;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1a: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_40 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_40 <= w_sys_tmp477;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h20: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_41 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_41 <= w_sys_tmp688;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h20: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_42 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_42 <= w_sys_tmp689;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h20: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_43 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_43 <= w_sys_tmp690;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h20: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_44 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_44 <= w_sys_tmp691;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h20: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_45 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_45 <= w_sys_tmp692;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_46 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_46 <= w_sys_tmp903;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_47 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_47 <= w_sys_tmp904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_48 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_48 <= w_sys_tmp905;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_49 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_49 <= w_sys_tmp906;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_50 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_50 <= w_sys_tmp907;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h31: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_51 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_51 <= w_sys_tmp1122;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h31: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_52 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_52 <= w_sys_tmp1123;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h31: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_53 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_53 <= w_sys_tmp1124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h31: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_54 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_54 <= w_sys_tmp1125;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h31: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_55 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_55 <= w_sys_tmp1126;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_56 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_56 <= w_sys_tmp1337;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_57 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_57 <= w_sys_tmp1338;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_58 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_58 <= w_sys_tmp1339;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_59 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_59 <= w_sys_tmp1340;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h37: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_60 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_60 <= w_sys_tmp1341;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_61 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_61 <= w_sys_tmp1552;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_62 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_62 <= w_sys_tmp1553;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_63 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_63 <= w_sys_tmp1554;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_64 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_64 <= w_sys_tmp1555;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_65 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_65 <= w_sys_tmp1556;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h43: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_66 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_66 <= w_sys_tmp1767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h43: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_67 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_67 <= w_sys_tmp1768;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h43: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_68 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_68 <= w_sys_tmp1769;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h43: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_69 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_69 <= w_sys_tmp1770;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h43: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_70 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_70 <= w_sys_tmp1771;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h57: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_71 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_run_copy0_j_71 <= w_sys_tmp2020;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h57: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_72 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_run_copy1_j_72 <= w_sys_tmp2021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h57: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_73 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_run_copy2_j_73 <= w_sys_tmp2022;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h5d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_74 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_run_copy0_j_74 <= w_sys_tmp2193;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h5d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_75 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_run_copy1_j_75 <= w_sys_tmp2194;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h5d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_76 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_run_copy2_j_76 <= w_sys_tmp2195;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h63: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_77 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_run_copy0_j_77 <= w_sys_tmp2366;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h63: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_78 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_run_copy1_j_78 <= w_sys_tmp2367;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h63: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_79 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_run_copy2_j_79 <= w_sys_tmp2368;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h69: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_80 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_run_copy0_j_80 <= w_sys_tmp2539;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h69: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_81 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_run_copy1_j_81 <= w_sys_tmp2540;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h69: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_82 <= r_run_j_13;

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_run_copy2_j_82 <= w_sys_tmp2541;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp896[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_datain <= w_sys_tmp899;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub03_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp888[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_V_datain <= w_sys_tmp891;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub03_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp880[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_datain <= w_sys_tmp883;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub03_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp1968[8:0] );

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2535[8:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2520[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub03_result_datain <= w_sys_tmp1970;

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub03_result_datain <= w_sys_tmp2524;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp681[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_datain <= w_sys_tmp684;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub02_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp673[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_V_datain <= w_sys_tmp676;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub02_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp665[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_datain <= w_sys_tmp668;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub02_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1990[8:0] );

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1980[8:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp1968[8:0] );

									end
								end

							endcase
						end

						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2362[8:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2347[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub02_result_datain <= w_sys_tmp2351;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'h2)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp466[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_datain <= w_sys_tmp469;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub01_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp458[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_V_datain <= w_sys_tmp461;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub01_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp450[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_datain <= w_sys_tmp453;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub01_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1985[8:0] );

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1990[8:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1974[8:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1980[8:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp1962[8:0] );

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2174[8:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2189[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub01_result_datain <= w_sys_tmp1976;

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'h7)) begin
										r_sub01_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sub01_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub01_result_datain <= w_sys_tmp2178;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h5<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp251[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_datain <= w_sys_tmp254;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub00_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp243[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_V_datain <= w_sys_tmp246;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub00_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp235[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_datain <= w_sys_tmp238;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub00_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1985[14:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1974[14:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1962[14:0] );

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2016[14:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2001[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_datain <= w_sys_tmp1964;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub00_result_datain <= w_sys_tmp2005;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h4)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h26)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h27)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp1760[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_datain <= w_sys_tmp1763;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub07_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1752[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_V_datain <= w_sys_tmp1755;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub07_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1744[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_datain <= w_sys_tmp1747;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub07_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2525[8:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2530[8:0] );

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2710[8:0] );

									end
									else
									if((r_sys_run_step==6'h4)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2722[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub07_result_datain <= w_sys_tmp2534;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub07_result_datain <= w_sys_tmp2712;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h6d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h4)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp1545[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_datain <= w_sys_tmp1548;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub06_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1537[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_V_datain <= w_sys_tmp1540;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub06_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1529[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_datain <= w_sys_tmp1532;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub06_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2357[8:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2352[8:0] );

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2710[8:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2722[8:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2705[8:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2716[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub06_result_datain <= w_sys_tmp2361;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub06_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub06_result_datain <= w_sys_tmp2695;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h67: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp1330[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_datain <= w_sys_tmp1333;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub05_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1322[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_V_datain <= w_sys_tmp1325;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub05_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1314[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_datain <= w_sys_tmp1317;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub05_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2179[8:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2184[8:0] );

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2699[8:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2705[8:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2716[8:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2693[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub05_result_datain <= w_sys_tmp2188;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub05_result_datain <= w_sys_tmp2701;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub05_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1115[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_datain <= w_sys_tmp1118;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub04_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1107[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_V_datain <= w_sys_tmp1110;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub04_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1099[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_datain <= w_sys_tmp1102;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub04_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2006[8:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2011[8:0] );

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2699[8:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2693[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub04_result_datain <= w_sys_tmp2015;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub04_result_datain <= w_sys_tmp2695;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h29)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h24)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h75: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h4)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						7'h73: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_tmp0_float <= w_sub07_result_dataout;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp1_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sys_tmp1_float <= w_sub00_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h19)) begin
										r_sys_tmp2_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h17)) begin
										r_sys_tmp3_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h19)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
