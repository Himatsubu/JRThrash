/*
TimeStamp:	2016/4/18		11:47
*/


module c1_unroll(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg  signed [31:0] r_ip_Multint_multiplicand_0;
	reg  signed [31:0] r_ip_Multint_multiplier_0;
	wire signed [63:0] w_ip_Multint_product_0;
	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_1;
	wire        [31:0] w_ip_FixedToFloat_floating_1;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_2;
	wire        [31:0] w_ip_FixedToFloat_floating_2;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_3;
	wire        [31:0] w_ip_FixedToFloat_floating_3;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_4;
	wire        [31:0] w_ip_FixedToFloat_floating_4;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_5;
	wire        [31:0] w_ip_FixedToFloat_floating_5;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_6;
	wire        [31:0] w_ip_FixedToFloat_floating_6;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_7;
	wire        [31:0] w_ip_FixedToFloat_floating_7;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_8;
	wire        [31:0] w_ip_FixedToFloat_floating_8;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_9;
	wire        [31:0] w_ip_FixedToFloat_floating_9;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 1:0] r_sys_run_stage;
	reg         [ 7:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 1:0] w_sys_run_stage_p1;
	wire        [ 7:0] w_sys_run_step_p1;
	wire signed [ 8:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [ 8:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [ 8:0] w_fld_uu_1_addr_0;
	wire        [31:0] w_fld_uu_1_datain_0;
	wire        [31:0] w_fld_uu_1_dataout_0;
	wire               w_fld_uu_1_r_w_0;
	wire               w_fld_uu_1_ce_0;
	reg  signed [ 8:0] r_fld_uu_1_addr_1;
	reg         [31:0] r_fld_uu_1_datain_1;
	wire        [31:0] w_fld_uu_1_dataout_1;
	reg                r_fld_uu_1_r_w_1;
	wire               w_fld_uu_1_ce_1;
	wire signed [ 8:0] w_fld_q_2_addr_0;
	wire        [31:0] w_fld_q_2_datain_0;
	wire        [31:0] w_fld_q_2_dataout_0;
	wire               w_fld_q_2_r_w_0;
	wire               w_fld_q_2_ce_0;
	reg  signed [ 8:0] r_fld_q_2_addr_1;
	reg         [31:0] r_fld_q_2_datain_1;
	wire        [31:0] w_fld_q_2_dataout_1;
	reg                r_fld_q_2_r_w_1;
	wire               w_fld_q_2_ce_1;
	reg  signed [31:0] r_run_k_3;
	reg  signed [31:0] r_run_j_4;
	reg  signed [31:0] r_run_n_5;
	reg  signed [31:0] r_run_mx_6;
	reg  signed [31:0] r_run_my_7;
	reg         [31:0] r_run_dt_8;
	reg         [31:0] r_run_dx_9;
	reg         [31:0] r_run_dy_10;
	reg         [31:0] r_run_r1_11;
	reg         [31:0] r_run_r2_12;
	reg  signed [31:0] r_run_kx_13;
	reg  signed [31:0] r_run_ky_14;
	reg  signed [31:0] r_run_nlast_15;
	reg  signed [31:0] r_run_copy0_j_16;
	reg  signed [31:0] r_run_copy1_j_17;
	reg  signed [31:0] r_run_copy2_j_18;
	reg  signed [31:0] r_run_copy0_j_19;
	reg  signed [31:0] r_run_copy0_j_20;
	reg  signed [31:0] r_run_copy1_j_21;
	reg  signed [31:0] r_run_copy2_j_22;
	reg  signed [31:0] r_run_copy3_j_23;
	reg  signed [31:0] r_run_copy4_j_24;
	reg  signed [31:0] r_run_copy5_j_25;
	reg  signed [31:0] r_run_copy6_j_26;
	reg  signed [31:0] r_run_copy7_j_27;
	reg  signed [31:0] r_run_copy0_j_28;
	reg  signed [31:0] r_sys_tmp0_int;
	reg  signed [31:0] r_sys_tmp1_int;
	reg  signed [31:0] r_sys_tmp2_int;
	reg  signed [31:0] r_sys_tmp3_int;
	reg  signed [31:0] r_sys_tmp4_int;
	reg  signed [31:0] r_sys_tmp5_int;
	reg  signed [31:0] r_sys_tmp6_int;
	reg  signed [31:0] r_sys_tmp7_int;
	reg  signed [31:0] r_sys_tmp8_int;
	reg  signed [31:0] r_sys_tmp9_int;
	reg  signed [31:0] r_sys_tmp10_int;
	reg  signed [31:0] r_sys_tmp11_int;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp9;
	wire               w_sys_tmp11;
	wire               w_sys_tmp12;
	wire signed [31:0] w_sys_tmp13;
	wire               w_sys_tmp14;
	wire               w_sys_tmp15;
	wire signed [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire        [31:0] w_sys_tmp20;
	wire        [31:0] w_sys_tmp21;
	wire        [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire signed [31:0] w_sys_tmp26;
	wire        [31:0] w_sys_tmp29;
	wire signed [31:0] w_sys_tmp35;
	wire signed [31:0] w_sys_tmp36;
	wire signed [31:0] w_sys_tmp37;
	wire signed [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp87;
	wire signed [31:0] w_sys_tmp88;
	wire               w_sys_tmp434;
	wire               w_sys_tmp435;
	wire signed [31:0] w_sys_tmp436;
	wire               w_sys_tmp437;
	wire               w_sys_tmp438;
	wire signed [31:0] w_sys_tmp441;
	wire signed [31:0] w_sys_tmp442;
	wire        [31:0] w_sys_tmp443;
	wire signed [31:0] w_sys_tmp445;
	wire signed [31:0] w_sys_tmp446;
	wire        [31:0] w_sys_tmp448;
	wire signed [31:0] w_sys_tmp449;
	wire               w_sys_tmp450;
	wire               w_sys_tmp451;
	wire signed [31:0] w_sys_tmp454;
	wire signed [31:0] w_sys_tmp455;
	wire signed [31:0] w_sys_tmp456;
	wire        [31:0] w_sys_tmp457;
	wire signed [31:0] w_sys_tmp459;
	wire        [31:0] w_sys_tmp462;
	wire signed [31:0] w_sys_tmp463;
	wire signed [31:0] w_sys_tmp464;
	wire signed [31:0] w_sys_tmp681;
	wire               w_sys_tmp682;
	wire               w_sys_tmp683;
	wire signed [31:0] w_sys_tmp684;
	wire signed [31:0] w_sys_tmp685;
	wire signed [31:0] w_sys_tmp686;
	wire               w_sys_tmp687;
	wire               w_sys_tmp688;
	wire signed [31:0] w_sys_tmp689;
	wire signed [31:0] w_sys_tmp692;
	wire signed [31:0] w_sys_tmp693;
	wire signed [31:0] w_sys_tmp694;
	wire        [31:0] w_sys_tmp695;
	wire        [31:0] w_sys_tmp699;
	wire signed [31:0] w_sys_tmp704;
	wire        [31:0] w_sys_tmp707;
	wire        [31:0] w_sys_tmp708;
	wire signed [31:0] w_sys_tmp714;
	wire signed [31:0] w_sys_tmp718;
	wire signed [31:0] w_sys_tmp728;
	wire        [31:0] w_sys_tmp733;
	wire signed [31:0] w_sys_tmp737;
	wire signed [31:0] w_sys_tmp738;
	wire signed [31:0] w_sys_tmp739;
	wire signed [31:0] w_sys_tmp740;
	wire signed [31:0] w_sys_tmp741;
	wire signed [31:0] w_sys_tmp742;
	wire signed [31:0] w_sys_tmp744;
	wire signed [31:0] w_sys_tmp745;
	wire signed [31:0] w_sys_tmp1705;
	wire               w_sys_tmp1706;
	wire               w_sys_tmp1707;
	wire signed [31:0] w_sys_tmp1708;
	wire signed [31:0] w_sys_tmp1709;
	wire signed [31:0] w_sys_tmp1710;
	wire               w_sys_tmp1711;
	wire               w_sys_tmp1712;
	wire signed [31:0] w_sys_tmp1713;
	wire signed [31:0] w_sys_tmp1716;
	wire signed [31:0] w_sys_tmp1717;
	wire signed [31:0] w_sys_tmp1718;
	wire        [31:0] w_sys_tmp1719;
	wire signed [31:0] w_sys_tmp1723;
	wire signed [31:0] w_sys_tmp1724;
	wire signed [31:0] w_sys_tmp1888;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 2'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 8'h1);
	assign w_fld_u_0_addr_0 = 9'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_fld_uu_1_addr_0 = 9'sh0;
	assign w_fld_uu_1_datain_0 = 32'h0;
	assign w_fld_uu_1_r_w_0 = 1'h0;
	assign w_fld_uu_1_ce_0 = w_sys_ce;
	assign w_fld_uu_1_ce_1 = w_sys_ce;
	assign w_fld_q_2_addr_0 = 9'sh0;
	assign w_fld_q_2_datain_0 = 32'h0;
	assign w_fld_q_2_r_w_0 = 1'h0;
	assign w_fld_q_2_ce_0 = w_sys_ce;
	assign w_fld_q_2_ce_1 = w_sys_ce;
	assign w_sys_tmp1 = 32'sh00000014;
	assign w_sys_tmp3 = 32'sh00000015;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'sh00000190;
	assign w_sys_tmp7 = 32'h3d4ccccd;
	assign w_sys_tmp9 = 32'h3e4ccccd;
	assign w_sys_tmp11 = ( !w_sys_tmp12 );
	assign w_sys_tmp12 = (r_run_my_7 < r_run_k_3);
	assign w_sys_tmp13 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp14 = ( !w_sys_tmp15 );
	assign w_sys_tmp15 = (r_run_mx_6 < r_run_j_4);
	assign w_sys_tmp18 = $signed( w_ip_Multint_product_0[31:0] );
	assign w_sys_tmp19 = 32'sh00000015;
	assign w_sys_tmp20 = w_ip_MultFloat_product_0;
	assign w_sys_tmp21 = 32'h42c80000;
	assign w_sys_tmp22 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp23 = (r_run_copy2_j_18 - w_sys_intOne);
	assign w_sys_tmp24 = (r_run_k_3 - w_sys_intOne);
	assign w_sys_tmp26 = (w_sys_tmp18 + r_run_k_3);
	assign w_sys_tmp29 = 32'h0;
	assign w_sys_tmp35 = (r_run_copy0_j_16 + w_sys_intOne);
	assign w_sys_tmp36 = (r_run_copy1_j_17 + w_sys_intOne);
	assign w_sys_tmp37 = (r_run_copy2_j_18 + w_sys_intOne);
	assign w_sys_tmp38 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp87 = (w_sys_tmp88 - w_sys_intOne);
	assign w_sys_tmp88 = w_sys_tmp37;
	assign w_sys_tmp434 = ( !w_sys_tmp435 );
	assign w_sys_tmp435 = (r_run_nlast_15 < r_run_n_5);
	assign w_sys_tmp436 = (r_run_n_5 + w_sys_intOne);
	assign w_sys_tmp437 = ( !w_sys_tmp438 );
	assign w_sys_tmp438 = (r_run_my_7 < r_run_k_3);
	assign w_sys_tmp441 = (w_sys_tmp442 + r_run_k_3);
	assign w_sys_tmp442 = 32'sh00000015;
	assign w_sys_tmp443 = 32'h3f000000;
	assign w_sys_tmp445 = (w_sys_tmp446 + r_run_k_3);
	assign w_sys_tmp446 = $signed( w_ip_Multint_product_0[31:0] );
	assign w_sys_tmp448 = 32'h0;
	assign w_sys_tmp449 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp450 = ( !w_sys_tmp451 );
	assign w_sys_tmp451 = (r_run_mx_6 < r_run_j_4);
	assign w_sys_tmp454 = (w_sys_tmp455 + w_sys_intOne);
	assign w_sys_tmp455 = $signed( w_ip_Multint_product_0[31:0] );
	assign w_sys_tmp456 = 32'sh00000015;
	assign w_sys_tmp457 = 32'h3f800000;
	assign w_sys_tmp459 = (w_sys_tmp455 + r_run_my_7);
	assign w_sys_tmp462 = 32'h0;
	assign w_sys_tmp463 = (r_run_copy0_j_19 + w_sys_intOne);
	assign w_sys_tmp464 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp681 = 32'sh00000002;
	assign w_sys_tmp682 = ( !w_sys_tmp683 );
	assign w_sys_tmp683 = (w_sys_tmp684 < r_run_k_3);
	assign w_sys_tmp684 = (r_run_my_7 - w_sys_intOne);
	assign w_sys_tmp685 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp686 = 32'sh00000002;
	assign w_sys_tmp687 = ( !w_sys_tmp688 );
	assign w_sys_tmp688 = (w_sys_tmp689 < r_run_j_4);
	assign w_sys_tmp689 = (r_run_mx_6 - w_sys_intOne);
	assign w_sys_tmp692 = (w_sys_tmp693 + r_run_k_3);
	assign w_sys_tmp693 = $signed( w_ip_Multint_product_0[31:0] );
	assign w_sys_tmp694 = 32'sh00000015;
	assign w_sys_tmp695 = w_ip_AddFloat_result_0;
	assign w_sys_tmp699 = w_ip_MultFloat_product_0;
	assign w_sys_tmp704 = (r_run_copy6_j_26 + w_sys_intOne);
	assign w_sys_tmp707 = 32'h40000000;
	assign w_sys_tmp708 = w_fld_u_0_dataout_1;
	assign w_sys_tmp714 = (r_run_copy4_j_24 - w_sys_intOne);
	assign w_sys_tmp718 = (w_sys_tmp692 + w_sys_intOne);
	assign w_sys_tmp728 = (w_sys_tmp692 - w_sys_intOne);
	assign w_sys_tmp733 = w_fld_q_2_dataout_1;
	assign w_sys_tmp737 = (r_run_copy0_j_20 + w_sys_intOne);
	assign w_sys_tmp738 = (r_run_copy1_j_21 + w_sys_intOne);
	assign w_sys_tmp739 = (r_run_copy2_j_22 + w_sys_intOne);
	assign w_sys_tmp740 = (r_run_copy3_j_23 + w_sys_intOne);
	assign w_sys_tmp741 = (r_run_copy4_j_24 + w_sys_intOne);
	assign w_sys_tmp742 = (r_run_copy5_j_25 + w_sys_intOne);
	assign w_sys_tmp744 = (r_run_copy7_j_27 + w_sys_intOne);
	assign w_sys_tmp745 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp1705 = 32'sh00000002;
	assign w_sys_tmp1706 = ( !w_sys_tmp1707 );
	assign w_sys_tmp1707 = (w_sys_tmp1708 < r_run_k_3);
	assign w_sys_tmp1708 = (r_run_my_7 - w_sys_intOne);
	assign w_sys_tmp1709 = (r_run_k_3 + w_sys_intOne);
	assign w_sys_tmp1710 = 32'sh00000002;
	assign w_sys_tmp1711 = ( !w_sys_tmp1712 );
	assign w_sys_tmp1712 = (w_sys_tmp1713 < r_run_j_4);
	assign w_sys_tmp1713 = (r_run_mx_6 - w_sys_intOne);
	assign w_sys_tmp1716 = (w_sys_tmp1717 + r_run_k_3);
	assign w_sys_tmp1717 = $signed( w_ip_Multint_product_0[31:0] );
	assign w_sys_tmp1718 = 32'sh00000015;
	assign w_sys_tmp1719 = w_fld_uu_1_dataout_1;
	assign w_sys_tmp1723 = (r_run_copy0_j_28 + w_sys_intOne);
	assign w_sys_tmp1724 = (r_run_j_4 + w_sys_intOne);
	assign w_sys_tmp1888 = (w_sys_tmp18 + r_run_k_3);


	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_uu_1(
			.clk (clock),
			.ce_0 (w_fld_uu_1_ce_0),
			.addr_0 (w_fld_uu_1_addr_0),
			.datain_0 (w_fld_uu_1_datain_0),
			.dataout_0 (w_fld_uu_1_dataout_0),
			.r_w_0 (w_fld_uu_1_r_w_0),
			.ce_1 (w_fld_uu_1_ce_1),
			.addr_1 (r_fld_uu_1_addr_1),
			.datain_1 (r_fld_uu_1_datain_1),
			.dataout_1 (w_fld_uu_1_dataout_1),
			.r_w_1 (r_fld_uu_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_q_2(
			.clk (clock),
			.ce_0 (w_fld_q_2_ce_0),
			.addr_0 (w_fld_q_2_addr_0),
			.datain_0 (w_fld_q_2_datain_0),
			.dataout_0 (w_fld_q_2_dataout_0),
			.r_w_0 (w_fld_q_2_r_w_0),
			.ce_1 (w_fld_q_2_ce_1),
			.addr_1 (r_fld_q_2_addr_1),
			.datain_1 (r_fld_q_2_datain_1),
			.dataout_1 (w_fld_q_2_dataout_1),
			.r_w_1 (r_fld_q_2_r_w_1)
		);

	Multint
		Multint_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_Multint_multiplicand_0),
			.b (r_ip_Multint_multiplier_0),
			.p (w_ip_Multint_product_0)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	FixedToFloat
		FixedToFloat_inst_1(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_1),
			.result (w_ip_FixedToFloat_floating_1)
		);

	FixedToFloat
		FixedToFloat_inst_2(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_2),
			.result (w_ip_FixedToFloat_floating_2)
		);

	FixedToFloat
		FixedToFloat_inst_3(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_3),
			.result (w_ip_FixedToFloat_floating_3)
		);

	FixedToFloat
		FixedToFloat_inst_4(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_4),
			.result (w_ip_FixedToFloat_floating_4)
		);

	FixedToFloat
		FixedToFloat_inst_5(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_5),
			.result (w_ip_FixedToFloat_floating_5)
		);

	FixedToFloat
		FixedToFloat_inst_6(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_6),
			.result (w_ip_FixedToFloat_floating_6)
		);

	FixedToFloat
		FixedToFloat_inst_7(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_7),
			.result (w_ip_FixedToFloat_floating_7)
		);

	FixedToFloat
		FixedToFloat_inst_8(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_8),
			.result (w_ip_FixedToFloat_floating_8)
		);

	FixedToFloat
		FixedToFloat_inst_9(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_9),
			.result (w_ip_FixedToFloat_floating_9)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h36)) begin
										r_ip_Multint_multiplicand_0 <= r_run_j_4;

									end
									else
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38)) begin
										r_ip_Multint_multiplicand_0 <= r_run_copy0_j_16;

									end
									else
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37)) begin
										r_ip_Multint_multiplicand_0 <= r_run_copy1_j_17;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_Multint_multiplicand_0 <= r_run_mx_6;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h2) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24)) begin
										r_ip_Multint_multiplicand_0 <= r_run_j_4;

									end
									else
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h25)) begin
										r_ip_Multint_multiplicand_0 <= r_run_copy0_j_19;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8f) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'h9d) || (8'h9f<=r_sys_run_step && r_sys_run_step<=8'haa)) begin
										r_ip_Multint_multiplicand_0 <= r_run_j_4;

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h87)) begin
										r_ip_Multint_multiplicand_0 <= r_run_copy1_j_21;

									end
									else
									if((r_sys_run_step==8'h4) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h70)) begin
										r_ip_Multint_multiplicand_0 <= r_run_copy5_j_25;

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h93)) begin
										r_ip_Multint_multiplicand_0 <= r_run_copy7_j_27;

									end
									else
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7d)) begin
										r_ip_Multint_multiplicand_0 <= w_sys_tmp714;

									end
									else
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h75)) begin
										r_ip_Multint_multiplicand_0 <= w_sys_tmp704;

									end
									else
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h74)) begin
										r_ip_Multint_multiplicand_0 <= r_run_copy2_j_22;

									end
									else
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7b)) begin
										r_ip_Multint_multiplicand_0 <= r_run_copy3_j_23;

									end
									else
									if((r_sys_run_step==8'h77) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'h9e)) begin
										r_ip_Multint_multiplicand_0 <= r_run_copy0_j_20;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h25)) begin
										r_ip_Multint_multiplicand_0 <= r_run_j_4;

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23)) begin
										r_ip_Multint_multiplicand_0 <= r_run_copy0_j_28;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h38)) begin
										r_ip_Multint_multiplier_0 <= w_sys_tmp19;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_ip_Multint_multiplier_0 <= w_sys_tmp442;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h25)) begin
										r_ip_Multint_multiplier_0 <= w_sys_tmp456;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'haa)) begin
										r_ip_Multint_multiplier_0 <= w_sys_tmp694;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h25)) begin
										r_ip_Multint_multiplier_0 <= w_sys_tmp1718;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h10) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h57)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h80)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h89) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'ha6)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'h8f)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h91) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'ha8)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'h83) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha4)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'h87) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'haa)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'h93)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h98)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h7c) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'h9a)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp708;

									end
									else
									if((r_sys_run_step==8'h25) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h84)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h86)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7f)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp695;

									end
									else
									if((r_sys_run_step==8'h8d) || (r_sys_run_step==8'ha0)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h33) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h9f)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'hd) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h8a)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h8b)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h95) || (r_sys_run_step==8'ha2)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'h2c) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h9d)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp14_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h15) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'h9d)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h19) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h70)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h1c) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h58)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp19_float[31], r_sys_tmp19_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'h9b)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h23) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h2b) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'h9f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h24) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'ha0) || (r_sys_run_step==8'ha1)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h84) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp708;

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp19_float[31], r_sys_tmp19_float[30:0] };

									end
									else
									if((r_sys_run_step==8'h31) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'h9e)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h2a) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h77)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'ha2) || (r_sys_run_step==8'ha4) || (r_sys_run_step==8'ha6) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'haa)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp699;

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp699[31], w_sys_tmp699[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h46)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==8'h14) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h41)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h24) || (r_sys_run_step==8'h32)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h49)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==8'h2c) || (r_sys_run_step==8'h38)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp34_float;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2a)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp21;

									end
									else
									if((r_sys_run_step==8'h1c) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3f)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4b)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h47)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h43)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==8'h20) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h3b)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==8'h28) || (r_sys_run_step==8'h35)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp26_float;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7b)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp707;

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h94)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r2_12;

									end
									else
									if((r_sys_run_step==8'h7e) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'ha5)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dt_8;

									end
									else
									if((r_sys_run_step==8'h1a) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h8a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r1_11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h33)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'h10) || (r_sys_run_step==8'h1f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'h11) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h45)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_dy_10;

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h8)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp22;

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h34)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp13_float;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2a)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_dx_9;

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h2b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp29_float;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h78)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h86)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp695;

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h94)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h90)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7b)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp708;

									end
									else
									if((r_sys_run_step==8'h7e) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'ha5)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp733;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h3<=r_sys_run_step && r_sys_run_step<=8'h11)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp87;

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1) || (r_sys_run_step==8'h2)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp23;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1) || (r_sys_run_step==8'h2)) begin
										r_ip_FixedToFloat_fixed_1 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_ip_FixedToFloat_fixed_2 <= w_sys_tmp87;

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1)) begin
										r_ip_FixedToFloat_fixed_2 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1)) begin
										r_ip_FixedToFloat_fixed_3 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1)) begin
										r_ip_FixedToFloat_fixed_4 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1)) begin
										r_ip_FixedToFloat_fixed_5 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1)) begin
										r_ip_FixedToFloat_fixed_6 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1)) begin
										r_ip_FixedToFloat_fixed_7 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1)) begin
										r_ip_FixedToFloat_fixed_8 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1)) begin
										r_ip_FixedToFloat_fixed_9 <= w_sys_tmp24;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h36: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp14) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h50)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp434) ? 6'h14 : 6'h36);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp437) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp450) ? 6'h1e : 6'h20);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2a)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp682) ? 6'h25 : 6'h2b);

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h26;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp687) ? 6'h29 : 6'h22);

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'haf)) begin
										r_sys_run_phase <= 6'h26;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h2c;

									end
								end

							endcase
						end

						6'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1706) ? 6'h30 : 6'h11);

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h2c;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h31;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1711) ? 6'h34 : 6'h2d);

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2a)) begin
										r_sys_run_phase <= 6'h31;

									end
								end

							endcase
						end

						6'h36: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h50)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2a)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'haf)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2a)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 8'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h4)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2a)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h29)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h26: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'haf)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'hae)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h2c: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h31: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h29)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h36: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp26[8:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp441[8:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp445[8:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp454[8:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp459[8:0] );

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp718[8:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (8'h8<=r_sys_run_step && r_sys_run_step<=8'hb) || (r_sys_run_step==8'hd) || (8'hf<=r_sys_run_step && r_sys_run_step<=8'h12) || (r_sys_run_step==8'h14) || (8'h16<=r_sys_run_step && r_sys_run_step<=8'h19) || (r_sys_run_step==8'h1b) || (8'h1d<=r_sys_run_step && r_sys_run_step<=8'h20) || (r_sys_run_step==8'h22) || (8'h24<=r_sys_run_step && r_sys_run_step<=8'h27) || (r_sys_run_step==8'h29) || (8'h2b<=r_sys_run_step && r_sys_run_step<=8'h2e) || (r_sys_run_step==8'h30) || (8'h32<=r_sys_run_step && r_sys_run_step<=8'h35) || (r_sys_run_step==8'h37) || (8'h39<=r_sys_run_step && r_sys_run_step<=8'h3c) || (r_sys_run_step==8'h3e) || (8'h40<=r_sys_run_step && r_sys_run_step<=8'h43) || (r_sys_run_step==8'h45) || (8'h47<=r_sys_run_step && r_sys_run_step<=8'h4a) || (r_sys_run_step==8'h4c) || (8'h4e<=r_sys_run_step && r_sys_run_step<=8'h51) || (r_sys_run_step==8'h53) || (8'h55<=r_sys_run_step && r_sys_run_step<=8'h58) || (r_sys_run_step==8'h5a) || (8'h5c<=r_sys_run_step && r_sys_run_step<=8'h5f) || (r_sys_run_step==8'h61) || (8'h63<=r_sys_run_step && r_sys_run_step<=8'h67) || (8'h69<=r_sys_run_step && r_sys_run_step<=8'h6c) || (8'h6e<=r_sys_run_step && r_sys_run_step<=8'h71) || (8'h73<=r_sys_run_step && r_sys_run_step<=8'h7b) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h98)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp692[8:0] );

									end
									else
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h8c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp728[8:0] );

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1716[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp29;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp443;

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp448;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp462;

									end
									else
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h29)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp457;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h2a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1719;

									end
									else
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h29)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp20_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h5)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h5<=r_sys_run_step && r_sys_run_step<=8'h2a)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h5<=r_sys_run_step && r_sys_run_step<=8'h7b) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h98)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2a)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h36: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3d)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp26[8:0] );

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h94) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha0) || (r_sys_run_step==8'ha2) || (8'ha4<=r_sys_run_step && r_sys_run_step<=8'haf)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp692[8:0] );

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h28)) begin
										r_fld_uu_1_addr_1 <= $signed( w_sys_tmp1716[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3d)) begin
										r_fld_uu_1_datain_1 <= w_sys_tmp29;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'haf)) begin
										r_fld_uu_1_datain_1 <= w_sys_tmp695;

									end
									else
									if((r_sys_run_step==8'haa)) begin
										r_fld_uu_1_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha7)) begin
										r_fld_uu_1_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'ha0) || (r_sys_run_step==8'ha8)) begin
										r_fld_uu_1_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'ha2)) begin
										r_fld_uu_1_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'h9a) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'had)) begin
										r_fld_uu_1_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'h97) || (r_sys_run_step==8'ha9) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'hae)) begin
										r_fld_uu_1_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'ha4)) begin
										r_fld_uu_1_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h9c) || (r_sys_run_step==8'ha6) || (r_sys_run_step==8'hab)) begin
										r_fld_uu_1_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h94)) begin
										r_fld_uu_1_datain_1 <= r_sys_tmp17_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_uu_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3d)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h94) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha0) || (r_sys_run_step==8'ha2) || (8'ha4<=r_sys_run_step && r_sys_run_step<=8'haf)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h28)) begin
										r_fld_uu_1_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_fld_uu_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_q_2_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h32) || (r_sys_run_step==8'h4d)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp8_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h3b) || (r_sys_run_step==8'h50)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp5_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp3_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp0_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp2_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h26) || (r_sys_run_step==8'h47)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp11_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp4_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h38) || (r_sys_run_step==8'h4f)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp6_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h35) || (r_sys_run_step==8'h4e)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp7_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h2a) || (r_sys_run_step==8'h4b)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp10_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp1_int[8:0] );

									end
									else
									if((r_sys_run_step==8'h2e) || (r_sys_run_step==8'h4c)) begin
										r_fld_q_2_addr_1 <= $signed( r_sys_tmp9_int[8:0] );

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'ha3)) begin
										r_fld_q_2_addr_1 <= $signed( w_sys_tmp692[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h26) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h49) || (8'h4b<=r_sys_run_step && r_sys_run_step<=8'h50)) begin
										r_fld_q_2_datain_1 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_q_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h26) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h49) || (8'h4b<=r_sys_run_step && r_sys_run_step<=8'h50)) begin
										r_fld_q_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'ha3)) begin
										r_fld_q_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h36: begin
							r_fld_q_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_3 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_3 <= w_sys_tmp13;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_3 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_run_k_3 <= w_sys_tmp449;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_3 <= w_sys_tmp681;

									end
								end

							endcase
						end

						6'h22: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_3 <= w_sys_tmp685;

									end
								end

							endcase
						end

						6'h2b: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_3 <= w_sys_tmp1705;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_3 <= w_sys_tmp1709;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h36)) begin
										r_run_j_4 <= w_sys_tmp38;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h2) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24)) begin
										r_run_j_4 <= w_sys_tmp464;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_4 <= w_sys_tmp686;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8f) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'h9d) || (8'h9f<=r_sys_run_step && r_sys_run_step<=8'haa)) begin
										r_run_j_4 <= w_sys_tmp745;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_4 <= w_sys_tmp1710;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h25)) begin
										r_run_j_4 <= w_sys_tmp1724;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_n_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_n_5 <= w_sys_tmp436;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_mx_6 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_my_7 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dt_8 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dx_9 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dy_10 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r1_11 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r2_12 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_kx_13 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_ky_14 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_nlast_15 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_16 <= r_run_j_4;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38)) begin
										r_run_copy0_j_16 <= w_sys_tmp35;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy1_j_17 <= r_run_j_4;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37)) begin
										r_run_copy1_j_17 <= w_sys_tmp36;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy2_j_18 <= r_run_j_4;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h12)) begin
										r_run_copy2_j_18 <= w_sys_tmp37;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1a: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_19 <= r_run_j_4;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h25)) begin
										r_run_copy0_j_19 <= w_sys_tmp463;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_20 <= r_run_j_4;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h77) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'h9e)) begin
										r_run_copy0_j_20 <= w_sys_tmp737;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy1_j_21 <= r_run_j_4;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h87)) begin
										r_run_copy1_j_21 <= w_sys_tmp738;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy2_j_22 <= r_run_j_4;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h74)) begin
										r_run_copy2_j_22 <= w_sys_tmp739;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy3_j_23 <= r_run_j_4;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7b)) begin
										r_run_copy3_j_23 <= w_sys_tmp740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy4_j_24 <= r_run_j_4;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7d)) begin
										r_run_copy4_j_24 <= w_sys_tmp741;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy5_j_25 <= r_run_j_4;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h4) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h70)) begin
										r_run_copy5_j_25 <= w_sys_tmp742;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy6_j_26 <= r_run_j_4;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h75)) begin
										r_run_copy6_j_26 <= w_sys_tmp704;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy7_j_27 <= r_run_j_4;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h93)) begin
										r_run_copy7_j_27 <= w_sys_tmp744;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h30: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_28 <= r_run_j_4;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h23)) begin
										r_run_copy0_j_28 <= w_sys_tmp1723;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h29)) begin
										r_sys_tmp0_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h23)) begin
										r_sys_tmp1_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_tmp2_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1d)) begin
										r_sys_tmp3_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sys_tmp4_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h3b)) begin
										r_sys_tmp5_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h14) || (r_sys_run_step==8'h38)) begin
										r_sys_tmp6_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h11) || (r_sys_run_step==8'h35)) begin
										r_sys_tmp7_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h32)) begin
										r_sys_tmp8_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hb) || (r_sys_run_step==8'h2f)) begin
										r_sys_tmp9_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'h2c)) begin
										r_sys_tmp10_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'h26)) begin
										r_sys_tmp11_int <= w_sys_tmp1888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sys_tmp0_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h68)) begin
										r_sys_tmp0_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h17)) begin
										r_sys_tmp1_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h75) || (r_sys_run_step==8'h78)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sys_tmp2_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6e) || (r_sys_run_step==8'h6f)) begin
										r_sys_tmp2_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_tmp3_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h61) || (r_sys_run_step==8'h9b)) begin
										r_sys_tmp3_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5a) || (r_sys_run_step==8'h98)) begin
										r_sys_tmp4_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h11)) begin
										r_sys_tmp5_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h53) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'ha3)) begin
										r_sys_tmp5_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hf)) begin
										r_sys_tmp6_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h4c) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'ha2)) begin
										r_sys_tmp6_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h9)) begin
										r_sys_tmp7_float <= w_ip_FixedToFloat_floating_1;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h45) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'ha0)) begin
										r_sys_tmp7_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp8_float <= w_ip_FixedToFloat_floating_9;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h37) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'ha6)) begin
										r_sys_tmp8_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp9_float <= w_ip_FixedToFloat_floating_1;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h30) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'hab)) begin
										r_sys_tmp9_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp10_float <= w_ip_FixedToFloat_floating_8;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3e) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'ha7)) begin
										r_sys_tmp10_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp11_float <= w_ip_FixedToFloat_floating_7;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h29) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9c) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha4) || (r_sys_run_step==8'ha9) || (r_sys_run_step==8'had)) begin
										r_sys_tmp11_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp12_float <= w_ip_FixedToFloat_floating_6;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h68)) begin
										r_sys_tmp12_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_sys_tmp12_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp13_float <= w_ip_FixedToFloat_floating_5;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h23) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h9d)) begin
										r_sys_tmp13_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp14_float <= w_ip_FixedToFloat_floating_2;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h11) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h61)) begin
										r_sys_tmp14_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==8'h76) || (r_sys_run_step==8'h77)) begin
										r_sys_tmp14_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp15_float <= w_ip_FixedToFloat_floating_4;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6b)) begin
										r_sys_tmp15_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7d)) begin
										r_sys_tmp15_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp16_float <= w_ip_FixedToFloat_floating_3;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8a) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h97)) begin
										r_sys_tmp16_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h70)) begin
										r_sys_tmp16_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp17_float <= w_ip_FixedToFloat_floating_1;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h65)) begin
										r_sys_tmp17_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==8'h71) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h88)) begin
										r_sys_tmp17_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp18_float <= w_ip_FixedToFloat_floating_3;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h9a)) begin
										r_sys_tmp18_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h72)) begin
										r_sys_tmp18_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==8'h80) || (r_sys_run_step==8'h81)) begin
										r_sys_tmp18_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp19_float <= w_ip_FixedToFloat_floating_9;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1c) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'ha0)) begin
										r_sys_tmp19_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp20_float <= w_ip_FixedToFloat_floating_8;

									end
								end

							endcase
						end

						6'h34: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h28)) begin
										r_sys_tmp20_float <= w_fld_uu_1_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp21_float <= w_ip_FixedToFloat_floating_7;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h81) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h98)) begin
										r_sys_tmp21_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h80)) begin
										r_sys_tmp21_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp22_float <= w_ip_FixedToFloat_floating_6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp23_float <= w_ip_FixedToFloat_floating_2;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp24_float <= w_ip_FixedToFloat_floating_5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp25_float <= w_ip_FixedToFloat_floating_4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1b) || (r_sys_run_step==8'h28)) begin
										r_sys_tmp26_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h24)) begin
										r_sys_tmp27_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hd) || (r_sys_run_step==8'h16)) begin
										r_sys_tmp28_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'h13)) begin
										r_sys_tmp29_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h15) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h30)) begin
										r_sys_tmp30_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h22)) begin
										r_sys_tmp31_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'hb) || (r_sys_run_step==8'h10)) begin
										r_sys_tmp31_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h36)) begin
										r_sys_tmp32_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hd) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h39)) begin
										r_sys_tmp33_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h2c)) begin
										r_sys_tmp34_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'he)) begin
										r_sys_tmp34_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hb) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h40)) begin
										r_sys_tmp35_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h3c)) begin
										r_sys_tmp36_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sys_tmp36_float <= w_ip_FixedToFloat_floating_2;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h42)) begin
										r_sys_tmp37_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h46)) begin
										r_sys_tmp38_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4a)) begin
										r_sys_tmp39_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
