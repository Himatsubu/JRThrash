/*
TimeStamp:	2016/10/20		16:0
*/


module P3_2dim(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 8:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [14:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [14:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [14:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [14:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [14:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [14:0] w_fld_V_3_addr_0;
	wire        [31:0] w_fld_V_3_datain_0;
	wire        [31:0] w_fld_V_3_dataout_0;
	wire               w_fld_V_3_r_w_0;
	wire               w_fld_V_3_ce_0;
	reg  signed [14:0] r_fld_V_3_addr_1;
	reg         [31:0] r_fld_V_3_datain_1;
	wire        [31:0] w_fld_V_3_dataout_1;
	reg                r_fld_V_3_r_w_1;
	wire               w_fld_V_3_ce_1;
	reg  signed [31:0] r_run_k_20;
	reg  signed [31:0] r_run_j_21;
	reg  signed [31:0] r_run_n_22;
	reg  signed [31:0] r_run_mx_23;
	reg  signed [31:0] r_run_my_24;
	reg         [31:0] r_run_dt_25;
	reg         [31:0] r_run_dx_26;
	reg         [31:0] r_run_dy_27;
	reg         [31:0] r_run_r1_28;
	reg         [31:0] r_run_r2_29;
	reg         [31:0] r_run_r3_30;
	reg         [31:0] r_run_r4_31;
	reg         [31:0] r_run_YY_32;
	reg  signed [31:0] r_run_kx_33;
	reg  signed [31:0] r_run_ky_34;
	reg  signed [31:0] r_run_nlast_35;
	reg  signed [31:0] r_run_tmpj_36;
	reg  signed [31:0] r_run_copy0_j_37;
	reg  signed [31:0] r_run_copy1_j_38;
	reg  signed [31:0] r_run_copy2_j_39;
	reg  signed [31:0] r_run_copy0_j_40;
	reg  signed [31:0] r_run_copy1_j_41;
	reg  signed [31:0] r_run_copy2_j_42;
	reg  signed [31:0] r_run_copy3_j_43;
	reg  signed [31:0] r_run_copy4_j_44;
	reg  signed [31:0] r_run_copy0_j_45;
	reg  signed [31:0] r_run_copy1_j_46;
	reg  signed [31:0] r_run_copy2_j_47;
	reg  signed [31:0] r_run_copy3_j_48;
	reg  signed [31:0] r_run_copy4_j_49;
	reg  signed [31:0] r_run_copy0_j_50;
	reg  signed [31:0] r_run_copy1_j_51;
	reg  signed [31:0] r_run_copy2_j_52;
	reg  signed [31:0] r_run_copy3_j_53;
	reg  signed [31:0] r_run_copy4_j_54;
	reg  signed [31:0] r_run_copy0_j_55;
	reg  signed [31:0] r_run_copy1_j_56;
	reg  signed [31:0] r_run_copy2_j_57;
	reg  signed [31:0] r_run_copy3_j_58;
	reg  signed [31:0] r_run_copy4_j_59;
	reg  signed [31:0] r_run_copy0_j_60;
	reg  signed [31:0] r_run_copy1_j_61;
	reg  signed [31:0] r_run_copy2_j_62;
	reg  signed [31:0] r_run_copy3_j_63;
	reg  signed [31:0] r_run_copy4_j_64;
	reg  signed [31:0] r_run_copy0_j_65;
	reg  signed [31:0] r_run_copy1_j_66;
	reg  signed [31:0] r_run_copy2_j_67;
	reg  signed [31:0] r_run_copy3_j_68;
	reg  signed [31:0] r_run_copy4_j_69;
	reg  signed [31:0] r_run_copy0_j_70;
	reg  signed [31:0] r_run_copy1_j_71;
	reg  signed [31:0] r_run_copy2_j_72;
	reg  signed [31:0] r_run_copy3_j_73;
	reg  signed [31:0] r_run_copy4_j_74;
	reg  signed [31:0] r_run_copy0_j_75;
	reg  signed [31:0] r_run_copy1_j_76;
	reg  signed [31:0] r_run_copy2_j_77;
	reg  signed [31:0] r_run_copy3_j_78;
	reg  signed [31:0] r_run_copy4_j_79;
	reg  signed [31:0] r_run_copy0_j_80;
	reg  signed [31:0] r_run_copy1_j_81;
	reg  signed [31:0] r_run_copy2_j_82;
	reg  signed [31:0] r_run_copy3_j_83;
	reg  signed [31:0] r_run_copy4_j_84;
	reg  signed [31:0] r_run_copy0_j_85;
	reg  signed [31:0] r_run_copy1_j_86;
	reg  signed [31:0] r_run_copy2_j_87;
	reg  signed [31:0] r_run_copy3_j_88;
	reg  signed [31:0] r_run_copy4_j_89;
	reg  signed [31:0] r_run_copy0_j_90;
	reg  signed [31:0] r_run_copy1_j_91;
	reg  signed [31:0] r_run_copy2_j_92;
	reg  signed [31:0] r_run_copy3_j_93;
	reg  signed [31:0] r_run_copy4_j_94;
	reg  signed [31:0] r_run_copy0_j_95;
	reg  signed [31:0] r_run_copy1_j_96;
	reg  signed [31:0] r_run_copy2_j_97;
	reg  signed [31:0] r_run_copy3_j_98;
	reg  signed [31:0] r_run_copy4_j_99;
	reg  signed [31:0] r_run_copy0_j_100;
	reg  signed [31:0] r_run_copy1_j_101;
	reg  signed [31:0] r_run_copy2_j_102;
	reg  signed [31:0] r_run_copy3_j_103;
	reg  signed [31:0] r_run_copy4_j_104;
	reg  signed [31:0] r_run_copy0_j_105;
	reg  signed [31:0] r_run_copy1_j_106;
	reg  signed [31:0] r_run_copy2_j_107;
	reg  signed [31:0] r_run_copy3_j_108;
	reg  signed [31:0] r_run_copy4_j_109;
	reg  signed [31:0] r_run_copy0_j_110;
	reg  signed [31:0] r_run_copy1_j_111;
	reg  signed [31:0] r_run_copy2_j_112;
	reg  signed [31:0] r_run_copy3_j_113;
	reg  signed [31:0] r_run_copy4_j_114;
	reg  signed [31:0] r_run_copy0_j_115;
	reg  signed [31:0] r_run_copy1_j_116;
	reg  signed [31:0] r_run_copy2_j_117;
	reg  signed [31:0] r_run_copy3_j_118;
	reg  signed [31:0] r_run_copy4_j_119;
	reg  signed [31:0] r_run_copy0_j_120;
	reg  signed [31:0] r_run_copy1_j_121;
	reg  signed [31:0] r_run_copy2_j_122;
	reg  signed [31:0] r_run_copy3_j_123;
	reg  signed [31:0] r_run_copy4_j_124;
	reg  signed [31:0] r_run_copy5_j_125;
	reg  signed [31:0] r_run_copy6_j_126;
	reg  signed [31:0] r_run_copy7_j_127;
	reg  signed [31:0] r_run_copy8_j_128;
	reg  signed [31:0] r_run_copy9_j_129;
	reg  signed [31:0] r_run_copy10_j_130;
	reg  signed [31:0] r_run_copy0_j_131;
	reg  signed [31:0] r_run_copy0_j_132;
	reg  signed [31:0] r_run_copy1_j_133;
	reg  signed [31:0] r_run_copy0_j_134;
	reg  signed [31:0] r_run_copy1_j_135;
	reg  signed [31:0] r_run_copy0_j_136;
	reg  signed [31:0] r_run_copy1_j_137;
	reg  signed [31:0] r_run_copy0_j_138;
	reg  signed [31:0] r_run_copy0_j_139;
	reg  signed [31:0] r_run_copy1_j_140;
	reg  signed [31:0] r_run_copy0_j_141;
	reg  signed [31:0] r_run_copy1_j_142;
	reg  signed [31:0] r_run_copy0_j_143;
	reg  signed [31:0] r_run_copy1_j_144;
	reg  signed [31:0] r_run_copy0_j_145;
	reg  signed [31:0] r_run_copy0_j_146;
	reg  signed [31:0] r_run_copy1_j_147;
	reg  signed [31:0] r_run_copy0_j_148;
	reg  signed [31:0] r_run_copy1_j_149;
	reg  signed [31:0] r_run_copy0_j_150;
	reg  signed [31:0] r_run_copy1_j_151;
	reg  signed [31:0] r_run_copy0_j_152;
	reg  signed [31:0] r_run_copy0_j_153;
	reg  signed [31:0] r_run_copy1_j_154;
	reg  signed [31:0] r_run_copy0_j_155;
	reg  signed [31:0] r_run_copy1_j_156;
	reg  signed [31:0] r_run_copy0_j_157;
	reg  signed [31:0] r_run_copy1_j_158;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [14:0] w_sub09_T_addr;
	reg  signed [14:0] r_sub09_T_addr;
	wire        [31:0] w_sub09_T_datain;
	reg         [31:0] r_sub09_T_datain;
	wire        [31:0] w_sub09_T_dataout;
	wire               w_sub09_T_r_w;
	reg                r_sub09_T_r_w;
	wire signed [14:0] w_sub09_V_addr;
	reg  signed [14:0] r_sub09_V_addr;
	wire        [31:0] w_sub09_V_datain;
	reg         [31:0] r_sub09_V_datain;
	wire        [31:0] w_sub09_V_dataout;
	wire               w_sub09_V_r_w;
	reg                r_sub09_V_r_w;
	wire signed [14:0] w_sub09_U_addr;
	reg  signed [14:0] r_sub09_U_addr;
	wire        [31:0] w_sub09_U_datain;
	reg         [31:0] r_sub09_U_datain;
	wire        [31:0] w_sub09_U_dataout;
	wire               w_sub09_U_r_w;
	reg                r_sub09_U_r_w;
	wire signed [14:0] w_sub09_result_addr;
	reg  signed [14:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [14:0] w_sub08_T_addr;
	reg  signed [14:0] r_sub08_T_addr;
	wire        [31:0] w_sub08_T_datain;
	reg         [31:0] r_sub08_T_datain;
	wire        [31:0] w_sub08_T_dataout;
	wire               w_sub08_T_r_w;
	reg                r_sub08_T_r_w;
	wire signed [14:0] w_sub08_V_addr;
	reg  signed [14:0] r_sub08_V_addr;
	wire        [31:0] w_sub08_V_datain;
	reg         [31:0] r_sub08_V_datain;
	wire        [31:0] w_sub08_V_dataout;
	wire               w_sub08_V_r_w;
	reg                r_sub08_V_r_w;
	wire signed [14:0] w_sub08_U_addr;
	reg  signed [14:0] r_sub08_U_addr;
	wire        [31:0] w_sub08_U_datain;
	reg         [31:0] r_sub08_U_datain;
	wire        [31:0] w_sub08_U_dataout;
	wire               w_sub08_U_r_w;
	reg                r_sub08_U_r_w;
	wire signed [14:0] w_sub08_result_addr;
	reg  signed [14:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [14:0] w_sub12_T_addr;
	reg  signed [14:0] r_sub12_T_addr;
	wire        [31:0] w_sub12_T_datain;
	reg         [31:0] r_sub12_T_datain;
	wire        [31:0] w_sub12_T_dataout;
	wire               w_sub12_T_r_w;
	reg                r_sub12_T_r_w;
	wire signed [14:0] w_sub12_V_addr;
	reg  signed [14:0] r_sub12_V_addr;
	wire        [31:0] w_sub12_V_datain;
	reg         [31:0] r_sub12_V_datain;
	wire        [31:0] w_sub12_V_dataout;
	wire               w_sub12_V_r_w;
	reg                r_sub12_V_r_w;
	wire signed [14:0] w_sub12_U_addr;
	reg  signed [14:0] r_sub12_U_addr;
	wire        [31:0] w_sub12_U_datain;
	reg         [31:0] r_sub12_U_datain;
	wire        [31:0] w_sub12_U_dataout;
	wire               w_sub12_U_r_w;
	reg                r_sub12_U_r_w;
	wire signed [14:0] w_sub12_result_addr;
	reg  signed [14:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [14:0] w_sub03_T_addr;
	reg  signed [14:0] r_sub03_T_addr;
	wire        [31:0] w_sub03_T_datain;
	reg         [31:0] r_sub03_T_datain;
	wire        [31:0] w_sub03_T_dataout;
	wire               w_sub03_T_r_w;
	reg                r_sub03_T_r_w;
	wire signed [14:0] w_sub03_V_addr;
	reg  signed [14:0] r_sub03_V_addr;
	wire        [31:0] w_sub03_V_datain;
	reg         [31:0] r_sub03_V_datain;
	wire        [31:0] w_sub03_V_dataout;
	wire               w_sub03_V_r_w;
	reg                r_sub03_V_r_w;
	wire signed [14:0] w_sub03_U_addr;
	reg  signed [14:0] r_sub03_U_addr;
	wire        [31:0] w_sub03_U_datain;
	reg         [31:0] r_sub03_U_datain;
	wire        [31:0] w_sub03_U_dataout;
	wire               w_sub03_U_r_w;
	reg                r_sub03_U_r_w;
	wire signed [14:0] w_sub03_result_addr;
	reg  signed [14:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [14:0] w_sub02_T_addr;
	reg  signed [14:0] r_sub02_T_addr;
	wire        [31:0] w_sub02_T_datain;
	reg         [31:0] r_sub02_T_datain;
	wire        [31:0] w_sub02_T_dataout;
	wire               w_sub02_T_r_w;
	reg                r_sub02_T_r_w;
	wire signed [14:0] w_sub02_V_addr;
	reg  signed [14:0] r_sub02_V_addr;
	wire        [31:0] w_sub02_V_datain;
	reg         [31:0] r_sub02_V_datain;
	wire        [31:0] w_sub02_V_dataout;
	wire               w_sub02_V_r_w;
	reg                r_sub02_V_r_w;
	wire signed [14:0] w_sub02_U_addr;
	reg  signed [14:0] r_sub02_U_addr;
	wire        [31:0] w_sub02_U_datain;
	reg         [31:0] r_sub02_U_datain;
	wire        [31:0] w_sub02_U_dataout;
	wire               w_sub02_U_r_w;
	reg                r_sub02_U_r_w;
	wire signed [14:0] w_sub02_result_addr;
	reg  signed [14:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [14:0] w_sub11_T_addr;
	reg  signed [14:0] r_sub11_T_addr;
	wire        [31:0] w_sub11_T_datain;
	reg         [31:0] r_sub11_T_datain;
	wire        [31:0] w_sub11_T_dataout;
	wire               w_sub11_T_r_w;
	reg                r_sub11_T_r_w;
	wire signed [14:0] w_sub11_V_addr;
	reg  signed [14:0] r_sub11_V_addr;
	wire        [31:0] w_sub11_V_datain;
	reg         [31:0] r_sub11_V_datain;
	wire        [31:0] w_sub11_V_dataout;
	wire               w_sub11_V_r_w;
	reg                r_sub11_V_r_w;
	wire signed [14:0] w_sub11_U_addr;
	reg  signed [14:0] r_sub11_U_addr;
	wire        [31:0] w_sub11_U_datain;
	reg         [31:0] r_sub11_U_datain;
	wire        [31:0] w_sub11_U_dataout;
	wire               w_sub11_U_r_w;
	reg                r_sub11_U_r_w;
	wire signed [14:0] w_sub11_result_addr;
	reg  signed [14:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [14:0] w_sub14_T_addr;
	reg  signed [14:0] r_sub14_T_addr;
	wire        [31:0] w_sub14_T_datain;
	reg         [31:0] r_sub14_T_datain;
	wire        [31:0] w_sub14_T_dataout;
	wire               w_sub14_T_r_w;
	reg                r_sub14_T_r_w;
	wire signed [14:0] w_sub14_V_addr;
	reg  signed [14:0] r_sub14_V_addr;
	wire        [31:0] w_sub14_V_datain;
	reg         [31:0] r_sub14_V_datain;
	wire        [31:0] w_sub14_V_dataout;
	wire               w_sub14_V_r_w;
	reg                r_sub14_V_r_w;
	wire signed [14:0] w_sub14_U_addr;
	reg  signed [14:0] r_sub14_U_addr;
	wire        [31:0] w_sub14_U_datain;
	reg         [31:0] r_sub14_U_datain;
	wire        [31:0] w_sub14_U_dataout;
	wire               w_sub14_U_r_w;
	reg                r_sub14_U_r_w;
	wire signed [14:0] w_sub14_result_addr;
	reg  signed [14:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [14:0] w_sub01_T_addr;
	reg  signed [14:0] r_sub01_T_addr;
	wire        [31:0] w_sub01_T_datain;
	reg         [31:0] r_sub01_T_datain;
	wire        [31:0] w_sub01_T_dataout;
	wire               w_sub01_T_r_w;
	reg                r_sub01_T_r_w;
	wire signed [14:0] w_sub01_V_addr;
	reg  signed [14:0] r_sub01_V_addr;
	wire        [31:0] w_sub01_V_datain;
	reg         [31:0] r_sub01_V_datain;
	wire        [31:0] w_sub01_V_dataout;
	wire               w_sub01_V_r_w;
	reg                r_sub01_V_r_w;
	wire signed [14:0] w_sub01_U_addr;
	reg  signed [14:0] r_sub01_U_addr;
	wire        [31:0] w_sub01_U_datain;
	reg         [31:0] r_sub01_U_datain;
	wire        [31:0] w_sub01_U_dataout;
	wire               w_sub01_U_r_w;
	reg                r_sub01_U_r_w;
	wire signed [14:0] w_sub01_result_addr;
	reg  signed [14:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [14:0] w_sub13_T_addr;
	reg  signed [14:0] r_sub13_T_addr;
	wire        [31:0] w_sub13_T_datain;
	reg         [31:0] r_sub13_T_datain;
	wire        [31:0] w_sub13_T_dataout;
	wire               w_sub13_T_r_w;
	reg                r_sub13_T_r_w;
	wire signed [14:0] w_sub13_V_addr;
	reg  signed [14:0] r_sub13_V_addr;
	wire        [31:0] w_sub13_V_datain;
	reg         [31:0] r_sub13_V_datain;
	wire        [31:0] w_sub13_V_dataout;
	wire               w_sub13_V_r_w;
	reg                r_sub13_V_r_w;
	wire signed [14:0] w_sub13_U_addr;
	reg  signed [14:0] r_sub13_U_addr;
	wire        [31:0] w_sub13_U_datain;
	reg         [31:0] r_sub13_U_datain;
	wire        [31:0] w_sub13_U_dataout;
	wire               w_sub13_U_r_w;
	reg                r_sub13_U_r_w;
	wire signed [14:0] w_sub13_result_addr;
	reg  signed [14:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [14:0] w_sub00_T_addr;
	reg  signed [14:0] r_sub00_T_addr;
	wire        [31:0] w_sub00_T_datain;
	reg         [31:0] r_sub00_T_datain;
	wire        [31:0] w_sub00_T_dataout;
	wire               w_sub00_T_r_w;
	reg                r_sub00_T_r_w;
	wire signed [14:0] w_sub00_V_addr;
	reg  signed [14:0] r_sub00_V_addr;
	wire        [31:0] w_sub00_V_datain;
	reg         [31:0] r_sub00_V_datain;
	wire        [31:0] w_sub00_V_dataout;
	wire               w_sub00_V_r_w;
	reg                r_sub00_V_r_w;
	wire signed [14:0] w_sub00_U_addr;
	reg  signed [14:0] r_sub00_U_addr;
	wire        [31:0] w_sub00_U_datain;
	reg         [31:0] r_sub00_U_datain;
	wire        [31:0] w_sub00_U_dataout;
	wire               w_sub00_U_r_w;
	reg                r_sub00_U_r_w;
	wire signed [14:0] w_sub00_result_addr;
	reg  signed [14:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [14:0] w_sub07_T_addr;
	reg  signed [14:0] r_sub07_T_addr;
	wire        [31:0] w_sub07_T_datain;
	reg         [31:0] r_sub07_T_datain;
	wire        [31:0] w_sub07_T_dataout;
	wire               w_sub07_T_r_w;
	reg                r_sub07_T_r_w;
	wire signed [14:0] w_sub07_V_addr;
	reg  signed [14:0] r_sub07_V_addr;
	wire        [31:0] w_sub07_V_datain;
	reg         [31:0] r_sub07_V_datain;
	wire        [31:0] w_sub07_V_dataout;
	wire               w_sub07_V_r_w;
	reg                r_sub07_V_r_w;
	wire signed [14:0] w_sub07_U_addr;
	reg  signed [14:0] r_sub07_U_addr;
	wire        [31:0] w_sub07_U_datain;
	reg         [31:0] r_sub07_U_datain;
	wire        [31:0] w_sub07_U_dataout;
	wire               w_sub07_U_r_w;
	reg                r_sub07_U_r_w;
	wire signed [14:0] w_sub07_result_addr;
	reg  signed [14:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [14:0] w_sub06_T_addr;
	reg  signed [14:0] r_sub06_T_addr;
	wire        [31:0] w_sub06_T_datain;
	reg         [31:0] r_sub06_T_datain;
	wire        [31:0] w_sub06_T_dataout;
	wire               w_sub06_T_r_w;
	reg                r_sub06_T_r_w;
	wire signed [14:0] w_sub06_V_addr;
	reg  signed [14:0] r_sub06_V_addr;
	wire        [31:0] w_sub06_V_datain;
	reg         [31:0] r_sub06_V_datain;
	wire        [31:0] w_sub06_V_dataout;
	wire               w_sub06_V_r_w;
	reg                r_sub06_V_r_w;
	wire signed [14:0] w_sub06_U_addr;
	reg  signed [14:0] r_sub06_U_addr;
	wire        [31:0] w_sub06_U_datain;
	reg         [31:0] r_sub06_U_datain;
	wire        [31:0] w_sub06_U_dataout;
	wire               w_sub06_U_r_w;
	reg                r_sub06_U_r_w;
	wire signed [14:0] w_sub06_result_addr;
	reg  signed [14:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [14:0] w_sub15_T_addr;
	reg  signed [14:0] r_sub15_T_addr;
	wire        [31:0] w_sub15_T_datain;
	reg         [31:0] r_sub15_T_datain;
	wire        [31:0] w_sub15_T_dataout;
	wire               w_sub15_T_r_w;
	reg                r_sub15_T_r_w;
	wire signed [14:0] w_sub15_V_addr;
	reg  signed [14:0] r_sub15_V_addr;
	wire        [31:0] w_sub15_V_datain;
	reg         [31:0] r_sub15_V_datain;
	wire        [31:0] w_sub15_V_dataout;
	wire               w_sub15_V_r_w;
	reg                r_sub15_V_r_w;
	wire signed [14:0] w_sub15_U_addr;
	reg  signed [14:0] r_sub15_U_addr;
	wire        [31:0] w_sub15_U_datain;
	reg         [31:0] r_sub15_U_datain;
	wire        [31:0] w_sub15_U_dataout;
	wire               w_sub15_U_r_w;
	reg                r_sub15_U_r_w;
	wire signed [14:0] w_sub15_result_addr;
	reg  signed [14:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [14:0] w_sub05_T_addr;
	reg  signed [14:0] r_sub05_T_addr;
	wire        [31:0] w_sub05_T_datain;
	reg         [31:0] r_sub05_T_datain;
	wire        [31:0] w_sub05_T_dataout;
	wire               w_sub05_T_r_w;
	reg                r_sub05_T_r_w;
	wire signed [14:0] w_sub05_V_addr;
	reg  signed [14:0] r_sub05_V_addr;
	wire        [31:0] w_sub05_V_datain;
	reg         [31:0] r_sub05_V_datain;
	wire        [31:0] w_sub05_V_dataout;
	wire               w_sub05_V_r_w;
	reg                r_sub05_V_r_w;
	wire signed [14:0] w_sub05_U_addr;
	reg  signed [14:0] r_sub05_U_addr;
	wire        [31:0] w_sub05_U_datain;
	reg         [31:0] r_sub05_U_datain;
	wire        [31:0] w_sub05_U_dataout;
	wire               w_sub05_U_r_w;
	reg                r_sub05_U_r_w;
	wire signed [14:0] w_sub05_result_addr;
	reg  signed [14:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [14:0] w_sub04_T_addr;
	reg  signed [14:0] r_sub04_T_addr;
	wire        [31:0] w_sub04_T_datain;
	reg         [31:0] r_sub04_T_datain;
	wire        [31:0] w_sub04_T_dataout;
	wire               w_sub04_T_r_w;
	reg                r_sub04_T_r_w;
	wire signed [14:0] w_sub04_V_addr;
	reg  signed [14:0] r_sub04_V_addr;
	wire        [31:0] w_sub04_V_datain;
	reg         [31:0] r_sub04_V_datain;
	wire        [31:0] w_sub04_V_dataout;
	wire               w_sub04_V_r_w;
	reg                r_sub04_V_r_w;
	wire signed [14:0] w_sub04_U_addr;
	reg  signed [14:0] r_sub04_U_addr;
	wire        [31:0] w_sub04_U_datain;
	reg         [31:0] r_sub04_U_datain;
	wire        [31:0] w_sub04_U_dataout;
	wire               w_sub04_U_r_w;
	reg                r_sub04_U_r_w;
	wire signed [14:0] w_sub04_result_addr;
	reg  signed [14:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [14:0] w_sub10_T_addr;
	reg  signed [14:0] r_sub10_T_addr;
	wire        [31:0] w_sub10_T_datain;
	reg         [31:0] r_sub10_T_datain;
	wire        [31:0] w_sub10_T_dataout;
	wire               w_sub10_T_r_w;
	reg                r_sub10_T_r_w;
	wire signed [14:0] w_sub10_V_addr;
	reg  signed [14:0] r_sub10_V_addr;
	wire        [31:0] w_sub10_V_datain;
	reg         [31:0] r_sub10_V_datain;
	wire        [31:0] w_sub10_V_dataout;
	wire               w_sub10_V_r_w;
	reg                r_sub10_V_r_w;
	wire signed [14:0] w_sub10_U_addr;
	reg  signed [14:0] r_sub10_U_addr;
	wire        [31:0] w_sub10_U_datain;
	reg         [31:0] r_sub10_U_datain;
	wire        [31:0] w_sub10_U_dataout;
	wire               w_sub10_U_r_w;
	reg                r_sub10_U_r_w;
	wire signed [14:0] w_sub10_result_addr;
	reg  signed [14:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire        [31:0] w_sys_tmp12;
	wire               w_sys_tmp13;
	wire               w_sys_tmp14;
	wire signed [31:0] w_sys_tmp15;
	wire               w_sys_tmp16;
	wire               w_sys_tmp17;
	wire        [31:0] w_sys_tmp19;
	wire        [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire signed [31:0] w_sys_tmp25;
	wire        [31:0] w_sys_tmp26;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp29;
	wire signed [31:0] w_sys_tmp33;
	wire signed [31:0] w_sys_tmp34;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire        [31:0] w_sys_tmp39;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp43;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire signed [31:0] w_sys_tmp49;
	wire        [31:0] w_sys_tmp129;
	wire               w_sys_tmp227;
	wire               w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire signed [31:0] w_sys_tmp230;
	wire               w_sys_tmp231;
	wire               w_sys_tmp232;
	wire signed [31:0] w_sys_tmp233;
	wire signed [31:0] w_sys_tmp236;
	wire signed [31:0] w_sys_tmp237;
	wire signed [31:0] w_sys_tmp238;
	wire        [31:0] w_sys_tmp239;
	wire signed [31:0] w_sys_tmp240;
	wire signed [31:0] w_sys_tmp241;
	wire signed [31:0] w_sys_tmp244;
	wire signed [31:0] w_sys_tmp245;
	wire        [31:0] w_sys_tmp247;
	wire signed [31:0] w_sys_tmp248;
	wire signed [31:0] w_sys_tmp249;
	wire signed [31:0] w_sys_tmp252;
	wire signed [31:0] w_sys_tmp253;
	wire        [31:0] w_sys_tmp255;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp257;
	wire signed [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp260;
	wire signed [31:0] w_sys_tmp261;
	wire signed [31:0] w_sys_tmp262;
	wire signed [31:0] w_sys_tmp263;
	wire signed [31:0] w_sys_tmp264;
	wire signed [31:0] w_sys_tmp445;
	wire               w_sys_tmp446;
	wire               w_sys_tmp447;
	wire signed [31:0] w_sys_tmp448;
	wire signed [31:0] w_sys_tmp451;
	wire signed [31:0] w_sys_tmp452;
	wire signed [31:0] w_sys_tmp453;
	wire        [31:0] w_sys_tmp454;
	wire signed [31:0] w_sys_tmp455;
	wire signed [31:0] w_sys_tmp456;
	wire signed [31:0] w_sys_tmp459;
	wire signed [31:0] w_sys_tmp460;
	wire        [31:0] w_sys_tmp462;
	wire signed [31:0] w_sys_tmp463;
	wire signed [31:0] w_sys_tmp464;
	wire signed [31:0] w_sys_tmp467;
	wire signed [31:0] w_sys_tmp468;
	wire        [31:0] w_sys_tmp470;
	wire signed [31:0] w_sys_tmp471;
	wire signed [31:0] w_sys_tmp472;
	wire signed [31:0] w_sys_tmp474;
	wire signed [31:0] w_sys_tmp475;
	wire signed [31:0] w_sys_tmp476;
	wire signed [31:0] w_sys_tmp477;
	wire signed [31:0] w_sys_tmp478;
	wire signed [31:0] w_sys_tmp479;
	wire signed [31:0] w_sys_tmp660;
	wire               w_sys_tmp661;
	wire               w_sys_tmp662;
	wire signed [31:0] w_sys_tmp663;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp667;
	wire signed [31:0] w_sys_tmp668;
	wire        [31:0] w_sys_tmp669;
	wire signed [31:0] w_sys_tmp670;
	wire signed [31:0] w_sys_tmp671;
	wire signed [31:0] w_sys_tmp674;
	wire signed [31:0] w_sys_tmp675;
	wire        [31:0] w_sys_tmp677;
	wire signed [31:0] w_sys_tmp678;
	wire signed [31:0] w_sys_tmp679;
	wire signed [31:0] w_sys_tmp682;
	wire signed [31:0] w_sys_tmp683;
	wire        [31:0] w_sys_tmp685;
	wire signed [31:0] w_sys_tmp686;
	wire signed [31:0] w_sys_tmp687;
	wire signed [31:0] w_sys_tmp689;
	wire signed [31:0] w_sys_tmp690;
	wire signed [31:0] w_sys_tmp691;
	wire signed [31:0] w_sys_tmp692;
	wire signed [31:0] w_sys_tmp693;
	wire signed [31:0] w_sys_tmp694;
	wire signed [31:0] w_sys_tmp875;
	wire               w_sys_tmp876;
	wire               w_sys_tmp877;
	wire signed [31:0] w_sys_tmp878;
	wire signed [31:0] w_sys_tmp881;
	wire signed [31:0] w_sys_tmp882;
	wire signed [31:0] w_sys_tmp883;
	wire        [31:0] w_sys_tmp884;
	wire signed [31:0] w_sys_tmp885;
	wire signed [31:0] w_sys_tmp886;
	wire signed [31:0] w_sys_tmp889;
	wire signed [31:0] w_sys_tmp890;
	wire        [31:0] w_sys_tmp892;
	wire signed [31:0] w_sys_tmp893;
	wire signed [31:0] w_sys_tmp894;
	wire signed [31:0] w_sys_tmp897;
	wire signed [31:0] w_sys_tmp898;
	wire        [31:0] w_sys_tmp900;
	wire signed [31:0] w_sys_tmp901;
	wire signed [31:0] w_sys_tmp902;
	wire signed [31:0] w_sys_tmp904;
	wire signed [31:0] w_sys_tmp905;
	wire signed [31:0] w_sys_tmp906;
	wire signed [31:0] w_sys_tmp907;
	wire signed [31:0] w_sys_tmp908;
	wire signed [31:0] w_sys_tmp909;
	wire signed [31:0] w_sys_tmp1090;
	wire               w_sys_tmp1091;
	wire               w_sys_tmp1092;
	wire signed [31:0] w_sys_tmp1093;
	wire signed [31:0] w_sys_tmp1094;
	wire               w_sys_tmp1095;
	wire               w_sys_tmp1096;
	wire signed [31:0] w_sys_tmp1097;
	wire signed [31:0] w_sys_tmp1100;
	wire signed [31:0] w_sys_tmp1101;
	wire signed [31:0] w_sys_tmp1102;
	wire        [31:0] w_sys_tmp1103;
	wire signed [31:0] w_sys_tmp1104;
	wire signed [31:0] w_sys_tmp1105;
	wire signed [31:0] w_sys_tmp1108;
	wire signed [31:0] w_sys_tmp1109;
	wire        [31:0] w_sys_tmp1111;
	wire signed [31:0] w_sys_tmp1112;
	wire signed [31:0] w_sys_tmp1113;
	wire signed [31:0] w_sys_tmp1116;
	wire signed [31:0] w_sys_tmp1117;
	wire        [31:0] w_sys_tmp1119;
	wire signed [31:0] w_sys_tmp1120;
	wire signed [31:0] w_sys_tmp1121;
	wire signed [31:0] w_sys_tmp1123;
	wire signed [31:0] w_sys_tmp1124;
	wire signed [31:0] w_sys_tmp1125;
	wire signed [31:0] w_sys_tmp1126;
	wire signed [31:0] w_sys_tmp1127;
	wire signed [31:0] w_sys_tmp1128;
	wire signed [31:0] w_sys_tmp1309;
	wire               w_sys_tmp1310;
	wire               w_sys_tmp1311;
	wire signed [31:0] w_sys_tmp1312;
	wire signed [31:0] w_sys_tmp1315;
	wire signed [31:0] w_sys_tmp1316;
	wire signed [31:0] w_sys_tmp1317;
	wire        [31:0] w_sys_tmp1318;
	wire signed [31:0] w_sys_tmp1319;
	wire signed [31:0] w_sys_tmp1320;
	wire signed [31:0] w_sys_tmp1323;
	wire signed [31:0] w_sys_tmp1324;
	wire        [31:0] w_sys_tmp1326;
	wire signed [31:0] w_sys_tmp1327;
	wire signed [31:0] w_sys_tmp1328;
	wire signed [31:0] w_sys_tmp1331;
	wire signed [31:0] w_sys_tmp1332;
	wire        [31:0] w_sys_tmp1334;
	wire signed [31:0] w_sys_tmp1335;
	wire signed [31:0] w_sys_tmp1336;
	wire signed [31:0] w_sys_tmp1338;
	wire signed [31:0] w_sys_tmp1339;
	wire signed [31:0] w_sys_tmp1340;
	wire signed [31:0] w_sys_tmp1341;
	wire signed [31:0] w_sys_tmp1342;
	wire signed [31:0] w_sys_tmp1343;
	wire signed [31:0] w_sys_tmp1524;
	wire               w_sys_tmp1525;
	wire               w_sys_tmp1526;
	wire signed [31:0] w_sys_tmp1527;
	wire signed [31:0] w_sys_tmp1530;
	wire signed [31:0] w_sys_tmp1531;
	wire signed [31:0] w_sys_tmp1532;
	wire        [31:0] w_sys_tmp1533;
	wire signed [31:0] w_sys_tmp1534;
	wire signed [31:0] w_sys_tmp1535;
	wire signed [31:0] w_sys_tmp1538;
	wire signed [31:0] w_sys_tmp1539;
	wire        [31:0] w_sys_tmp1541;
	wire signed [31:0] w_sys_tmp1542;
	wire signed [31:0] w_sys_tmp1543;
	wire signed [31:0] w_sys_tmp1546;
	wire signed [31:0] w_sys_tmp1547;
	wire        [31:0] w_sys_tmp1549;
	wire signed [31:0] w_sys_tmp1550;
	wire signed [31:0] w_sys_tmp1551;
	wire signed [31:0] w_sys_tmp1553;
	wire signed [31:0] w_sys_tmp1554;
	wire signed [31:0] w_sys_tmp1555;
	wire signed [31:0] w_sys_tmp1556;
	wire signed [31:0] w_sys_tmp1557;
	wire signed [31:0] w_sys_tmp1558;
	wire signed [31:0] w_sys_tmp1739;
	wire               w_sys_tmp1740;
	wire               w_sys_tmp1741;
	wire signed [31:0] w_sys_tmp1742;
	wire signed [31:0] w_sys_tmp1745;
	wire signed [31:0] w_sys_tmp1746;
	wire signed [31:0] w_sys_tmp1747;
	wire        [31:0] w_sys_tmp1748;
	wire signed [31:0] w_sys_tmp1749;
	wire signed [31:0] w_sys_tmp1750;
	wire signed [31:0] w_sys_tmp1753;
	wire signed [31:0] w_sys_tmp1754;
	wire        [31:0] w_sys_tmp1756;
	wire signed [31:0] w_sys_tmp1757;
	wire signed [31:0] w_sys_tmp1758;
	wire signed [31:0] w_sys_tmp1761;
	wire signed [31:0] w_sys_tmp1762;
	wire        [31:0] w_sys_tmp1764;
	wire signed [31:0] w_sys_tmp1765;
	wire signed [31:0] w_sys_tmp1766;
	wire signed [31:0] w_sys_tmp1768;
	wire signed [31:0] w_sys_tmp1769;
	wire signed [31:0] w_sys_tmp1770;
	wire signed [31:0] w_sys_tmp1771;
	wire signed [31:0] w_sys_tmp1772;
	wire signed [31:0] w_sys_tmp1773;
	wire signed [31:0] w_sys_tmp1954;
	wire               w_sys_tmp1955;
	wire               w_sys_tmp1956;
	wire signed [31:0] w_sys_tmp1957;
	wire signed [31:0] w_sys_tmp1958;
	wire               w_sys_tmp1959;
	wire               w_sys_tmp1960;
	wire signed [31:0] w_sys_tmp1961;
	wire signed [31:0] w_sys_tmp1964;
	wire signed [31:0] w_sys_tmp1965;
	wire signed [31:0] w_sys_tmp1966;
	wire        [31:0] w_sys_tmp1967;
	wire signed [31:0] w_sys_tmp1968;
	wire signed [31:0] w_sys_tmp1969;
	wire signed [31:0] w_sys_tmp1972;
	wire signed [31:0] w_sys_tmp1973;
	wire        [31:0] w_sys_tmp1975;
	wire signed [31:0] w_sys_tmp1976;
	wire signed [31:0] w_sys_tmp1977;
	wire signed [31:0] w_sys_tmp1980;
	wire signed [31:0] w_sys_tmp1981;
	wire        [31:0] w_sys_tmp1983;
	wire signed [31:0] w_sys_tmp1984;
	wire signed [31:0] w_sys_tmp1985;
	wire signed [31:0] w_sys_tmp1987;
	wire signed [31:0] w_sys_tmp1988;
	wire signed [31:0] w_sys_tmp1989;
	wire signed [31:0] w_sys_tmp1990;
	wire signed [31:0] w_sys_tmp1991;
	wire signed [31:0] w_sys_tmp1992;
	wire signed [31:0] w_sys_tmp2173;
	wire               w_sys_tmp2174;
	wire               w_sys_tmp2175;
	wire signed [31:0] w_sys_tmp2176;
	wire signed [31:0] w_sys_tmp2179;
	wire signed [31:0] w_sys_tmp2180;
	wire signed [31:0] w_sys_tmp2181;
	wire        [31:0] w_sys_tmp2182;
	wire signed [31:0] w_sys_tmp2183;
	wire signed [31:0] w_sys_tmp2184;
	wire signed [31:0] w_sys_tmp2187;
	wire signed [31:0] w_sys_tmp2188;
	wire        [31:0] w_sys_tmp2190;
	wire signed [31:0] w_sys_tmp2191;
	wire signed [31:0] w_sys_tmp2192;
	wire signed [31:0] w_sys_tmp2195;
	wire signed [31:0] w_sys_tmp2196;
	wire        [31:0] w_sys_tmp2198;
	wire signed [31:0] w_sys_tmp2199;
	wire signed [31:0] w_sys_tmp2200;
	wire signed [31:0] w_sys_tmp2202;
	wire signed [31:0] w_sys_tmp2203;
	wire signed [31:0] w_sys_tmp2204;
	wire signed [31:0] w_sys_tmp2205;
	wire signed [31:0] w_sys_tmp2206;
	wire signed [31:0] w_sys_tmp2207;
	wire signed [31:0] w_sys_tmp2388;
	wire               w_sys_tmp2389;
	wire               w_sys_tmp2390;
	wire signed [31:0] w_sys_tmp2391;
	wire signed [31:0] w_sys_tmp2394;
	wire signed [31:0] w_sys_tmp2395;
	wire signed [31:0] w_sys_tmp2396;
	wire        [31:0] w_sys_tmp2397;
	wire signed [31:0] w_sys_tmp2398;
	wire signed [31:0] w_sys_tmp2399;
	wire signed [31:0] w_sys_tmp2402;
	wire signed [31:0] w_sys_tmp2403;
	wire        [31:0] w_sys_tmp2405;
	wire signed [31:0] w_sys_tmp2406;
	wire signed [31:0] w_sys_tmp2407;
	wire signed [31:0] w_sys_tmp2410;
	wire signed [31:0] w_sys_tmp2411;
	wire        [31:0] w_sys_tmp2413;
	wire signed [31:0] w_sys_tmp2414;
	wire signed [31:0] w_sys_tmp2415;
	wire signed [31:0] w_sys_tmp2417;
	wire signed [31:0] w_sys_tmp2418;
	wire signed [31:0] w_sys_tmp2419;
	wire signed [31:0] w_sys_tmp2420;
	wire signed [31:0] w_sys_tmp2421;
	wire signed [31:0] w_sys_tmp2422;
	wire signed [31:0] w_sys_tmp2603;
	wire               w_sys_tmp2604;
	wire               w_sys_tmp2605;
	wire signed [31:0] w_sys_tmp2606;
	wire signed [31:0] w_sys_tmp2609;
	wire signed [31:0] w_sys_tmp2610;
	wire signed [31:0] w_sys_tmp2611;
	wire        [31:0] w_sys_tmp2612;
	wire signed [31:0] w_sys_tmp2613;
	wire signed [31:0] w_sys_tmp2614;
	wire signed [31:0] w_sys_tmp2617;
	wire signed [31:0] w_sys_tmp2618;
	wire        [31:0] w_sys_tmp2620;
	wire signed [31:0] w_sys_tmp2621;
	wire signed [31:0] w_sys_tmp2622;
	wire signed [31:0] w_sys_tmp2625;
	wire signed [31:0] w_sys_tmp2626;
	wire        [31:0] w_sys_tmp2628;
	wire signed [31:0] w_sys_tmp2629;
	wire signed [31:0] w_sys_tmp2630;
	wire signed [31:0] w_sys_tmp2632;
	wire signed [31:0] w_sys_tmp2633;
	wire signed [31:0] w_sys_tmp2634;
	wire signed [31:0] w_sys_tmp2635;
	wire signed [31:0] w_sys_tmp2636;
	wire signed [31:0] w_sys_tmp2637;
	wire signed [31:0] w_sys_tmp2818;
	wire               w_sys_tmp2819;
	wire               w_sys_tmp2820;
	wire signed [31:0] w_sys_tmp2821;
	wire signed [31:0] w_sys_tmp2822;
	wire               w_sys_tmp2823;
	wire               w_sys_tmp2824;
	wire signed [31:0] w_sys_tmp2825;
	wire signed [31:0] w_sys_tmp2828;
	wire signed [31:0] w_sys_tmp2829;
	wire signed [31:0] w_sys_tmp2830;
	wire        [31:0] w_sys_tmp2831;
	wire signed [31:0] w_sys_tmp2832;
	wire signed [31:0] w_sys_tmp2833;
	wire signed [31:0] w_sys_tmp2836;
	wire signed [31:0] w_sys_tmp2837;
	wire        [31:0] w_sys_tmp2839;
	wire signed [31:0] w_sys_tmp2840;
	wire signed [31:0] w_sys_tmp2841;
	wire signed [31:0] w_sys_tmp2844;
	wire signed [31:0] w_sys_tmp2845;
	wire        [31:0] w_sys_tmp2847;
	wire signed [31:0] w_sys_tmp2848;
	wire signed [31:0] w_sys_tmp2849;
	wire signed [31:0] w_sys_tmp2851;
	wire signed [31:0] w_sys_tmp2852;
	wire signed [31:0] w_sys_tmp2853;
	wire signed [31:0] w_sys_tmp2854;
	wire signed [31:0] w_sys_tmp2855;
	wire signed [31:0] w_sys_tmp2856;
	wire signed [31:0] w_sys_tmp3037;
	wire               w_sys_tmp3038;
	wire               w_sys_tmp3039;
	wire signed [31:0] w_sys_tmp3040;
	wire signed [31:0] w_sys_tmp3043;
	wire signed [31:0] w_sys_tmp3044;
	wire signed [31:0] w_sys_tmp3045;
	wire        [31:0] w_sys_tmp3046;
	wire signed [31:0] w_sys_tmp3047;
	wire signed [31:0] w_sys_tmp3048;
	wire signed [31:0] w_sys_tmp3051;
	wire signed [31:0] w_sys_tmp3052;
	wire        [31:0] w_sys_tmp3054;
	wire signed [31:0] w_sys_tmp3055;
	wire signed [31:0] w_sys_tmp3056;
	wire signed [31:0] w_sys_tmp3059;
	wire signed [31:0] w_sys_tmp3060;
	wire        [31:0] w_sys_tmp3062;
	wire signed [31:0] w_sys_tmp3063;
	wire signed [31:0] w_sys_tmp3064;
	wire signed [31:0] w_sys_tmp3066;
	wire signed [31:0] w_sys_tmp3067;
	wire signed [31:0] w_sys_tmp3068;
	wire signed [31:0] w_sys_tmp3069;
	wire signed [31:0] w_sys_tmp3070;
	wire signed [31:0] w_sys_tmp3071;
	wire signed [31:0] w_sys_tmp3252;
	wire               w_sys_tmp3253;
	wire               w_sys_tmp3254;
	wire signed [31:0] w_sys_tmp3255;
	wire signed [31:0] w_sys_tmp3258;
	wire signed [31:0] w_sys_tmp3259;
	wire signed [31:0] w_sys_tmp3260;
	wire        [31:0] w_sys_tmp3261;
	wire signed [31:0] w_sys_tmp3262;
	wire signed [31:0] w_sys_tmp3263;
	wire signed [31:0] w_sys_tmp3266;
	wire signed [31:0] w_sys_tmp3267;
	wire        [31:0] w_sys_tmp3269;
	wire signed [31:0] w_sys_tmp3270;
	wire signed [31:0] w_sys_tmp3271;
	wire signed [31:0] w_sys_tmp3274;
	wire signed [31:0] w_sys_tmp3275;
	wire        [31:0] w_sys_tmp3277;
	wire signed [31:0] w_sys_tmp3278;
	wire signed [31:0] w_sys_tmp3279;
	wire signed [31:0] w_sys_tmp3281;
	wire signed [31:0] w_sys_tmp3282;
	wire signed [31:0] w_sys_tmp3283;
	wire signed [31:0] w_sys_tmp3284;
	wire signed [31:0] w_sys_tmp3285;
	wire signed [31:0] w_sys_tmp3286;
	wire signed [31:0] w_sys_tmp3467;
	wire               w_sys_tmp3468;
	wire               w_sys_tmp3469;
	wire signed [31:0] w_sys_tmp3470;
	wire signed [31:0] w_sys_tmp3473;
	wire signed [31:0] w_sys_tmp3474;
	wire signed [31:0] w_sys_tmp3475;
	wire        [31:0] w_sys_tmp3476;
	wire signed [31:0] w_sys_tmp3477;
	wire signed [31:0] w_sys_tmp3478;
	wire signed [31:0] w_sys_tmp3481;
	wire signed [31:0] w_sys_tmp3482;
	wire        [31:0] w_sys_tmp3484;
	wire signed [31:0] w_sys_tmp3485;
	wire signed [31:0] w_sys_tmp3486;
	wire signed [31:0] w_sys_tmp3489;
	wire signed [31:0] w_sys_tmp3490;
	wire        [31:0] w_sys_tmp3492;
	wire signed [31:0] w_sys_tmp3493;
	wire signed [31:0] w_sys_tmp3494;
	wire signed [31:0] w_sys_tmp3496;
	wire signed [31:0] w_sys_tmp3497;
	wire signed [31:0] w_sys_tmp3498;
	wire signed [31:0] w_sys_tmp3499;
	wire signed [31:0] w_sys_tmp3500;
	wire signed [31:0] w_sys_tmp3501;
	wire               w_sys_tmp3682;
	wire               w_sys_tmp3683;
	wire signed [31:0] w_sys_tmp3684;
	wire signed [31:0] w_sys_tmp3685;
	wire               w_sys_tmp3686;
	wire               w_sys_tmp3687;
	wire signed [31:0] w_sys_tmp3688;
	wire signed [31:0] w_sys_tmp3691;
	wire signed [31:0] w_sys_tmp3692;
	wire        [31:0] w_sys_tmp3693;
	wire signed [31:0] w_sys_tmp3694;
	wire signed [31:0] w_sys_tmp3695;
	wire signed [31:0] w_sys_tmp3697;
	wire signed [31:0] w_sys_tmp3698;
	wire        [31:0] w_sys_tmp3699;
	wire signed [31:0] w_sys_tmp3700;
	wire signed [31:0] w_sys_tmp3701;
	wire signed [31:0] w_sys_tmp3703;
	wire signed [31:0] w_sys_tmp3704;
	wire        [31:0] w_sys_tmp3721;
	wire signed [31:0] w_sys_tmp3724;
	wire signed [31:0] w_sys_tmp3725;
	wire               w_sys_tmp3726;
	wire               w_sys_tmp3727;
	wire signed [31:0] w_sys_tmp3728;
	wire signed [31:0] w_sys_tmp3731;
	wire signed [31:0] w_sys_tmp3732;
	wire        [31:0] w_sys_tmp3733;
	wire signed [31:0] w_sys_tmp3734;
	wire signed [31:0] w_sys_tmp3735;
	wire signed [31:0] w_sys_tmp3737;
	wire signed [31:0] w_sys_tmp3738;
	wire        [31:0] w_sys_tmp3739;
	wire signed [31:0] w_sys_tmp3740;
	wire signed [31:0] w_sys_tmp3741;
	wire signed [31:0] w_sys_tmp3743;
	wire signed [31:0] w_sys_tmp3744;
	wire        [31:0] w_sys_tmp3761;
	wire signed [31:0] w_sys_tmp3764;
	wire signed [31:0] w_sys_tmp3765;
	wire               w_sys_tmp3766;
	wire               w_sys_tmp3767;
	wire signed [31:0] w_sys_tmp3768;
	wire signed [31:0] w_sys_tmp3771;
	wire signed [31:0] w_sys_tmp3772;
	wire        [31:0] w_sys_tmp3773;
	wire signed [31:0] w_sys_tmp3774;
	wire signed [31:0] w_sys_tmp3775;
	wire signed [31:0] w_sys_tmp3777;
	wire signed [31:0] w_sys_tmp3778;
	wire        [31:0] w_sys_tmp3779;
	wire signed [31:0] w_sys_tmp3780;
	wire signed [31:0] w_sys_tmp3781;
	wire signed [31:0] w_sys_tmp3783;
	wire signed [31:0] w_sys_tmp3784;
	wire        [31:0] w_sys_tmp3801;
	wire signed [31:0] w_sys_tmp3804;
	wire signed [31:0] w_sys_tmp3805;
	wire               w_sys_tmp3806;
	wire               w_sys_tmp3807;
	wire signed [31:0] w_sys_tmp3808;
	wire signed [31:0] w_sys_tmp3811;
	wire signed [31:0] w_sys_tmp3812;
	wire        [31:0] w_sys_tmp3813;
	wire signed [31:0] w_sys_tmp3814;
	wire signed [31:0] w_sys_tmp3815;
	wire signed [31:0] w_sys_tmp3817;
	wire signed [31:0] w_sys_tmp3818;
	wire        [31:0] w_sys_tmp3819;
	wire signed [31:0] w_sys_tmp3820;
	wire signed [31:0] w_sys_tmp3821;
	wire signed [31:0] w_sys_tmp3823;
	wire signed [31:0] w_sys_tmp3824;
	wire        [31:0] w_sys_tmp3841;
	wire signed [31:0] w_sys_tmp3842;
	wire signed [31:0] w_sys_tmp3843;
	wire signed [31:0] w_sys_tmp3844;
	wire signed [31:0] w_sys_tmp3845;
	wire               w_sys_tmp3846;
	wire               w_sys_tmp3847;
	wire signed [31:0] w_sys_tmp3848;
	wire signed [31:0] w_sys_tmp3851;
	wire signed [31:0] w_sys_tmp3852;
	wire signed [31:0] w_sys_tmp3853;
	wire signed [31:0] w_sys_tmp3854;
	wire        [31:0] w_sys_tmp3855;
	wire signed [31:0] w_sys_tmp3856;
	wire signed [31:0] w_sys_tmp3857;
	wire signed [31:0] w_sys_tmp3861;
	wire signed [31:0] w_sys_tmp3862;
	wire signed [31:0] w_sys_tmp3864;
	wire        [31:0] w_sys_tmp3865;
	wire signed [31:0] w_sys_tmp3866;
	wire signed [31:0] w_sys_tmp3867;
	wire signed [31:0] w_sys_tmp3871;
	wire signed [31:0] w_sys_tmp3872;
	wire signed [31:0] w_sys_tmp3874;
	wire signed [31:0] w_sys_tmp3875;
	wire signed [31:0] w_sys_tmp3876;
	wire signed [31:0] w_sys_tmp3880;
	wire signed [31:0] w_sys_tmp3881;
	wire signed [31:0] w_sys_tmp3883;
	wire signed [31:0] w_sys_tmp3885;
	wire signed [31:0] w_sys_tmp3886;
	wire signed [31:0] w_sys_tmp3890;
	wire signed [31:0] w_sys_tmp3891;
	wire signed [31:0] w_sys_tmp3893;
	wire signed [31:0] w_sys_tmp3894;
	wire signed [31:0] w_sys_tmp3895;
	wire signed [31:0] w_sys_tmp3899;
	wire signed [31:0] w_sys_tmp3900;
	wire signed [31:0] w_sys_tmp3902;
	wire        [31:0] w_sys_tmp3903;
	wire signed [31:0] w_sys_tmp3904;
	wire signed [31:0] w_sys_tmp3905;
	wire signed [31:0] w_sys_tmp3908;
	wire signed [31:0] w_sys_tmp3909;
	wire signed [31:0] w_sys_tmp3910;
	wire signed [31:0] w_sys_tmp3911;
	wire signed [31:0] w_sys_tmp3912;
	wire signed [31:0] w_sys_tmp3913;
	wire signed [31:0] w_sys_tmp3914;
	wire signed [31:0] w_sys_tmp3915;
	wire signed [31:0] w_sys_tmp3916;
	wire signed [31:0] w_sys_tmp3917;
	wire signed [31:0] w_sys_tmp3918;
	wire signed [31:0] w_sys_tmp3919;
	wire signed [31:0] w_sys_tmp4346;
	wire               w_sys_tmp4347;
	wire               w_sys_tmp4348;
	wire signed [31:0] w_sys_tmp4349;
	wire signed [31:0] w_sys_tmp4351;
	wire signed [31:0] w_sys_tmp4352;
	wire signed [31:0] w_sys_tmp4354;
	wire signed [31:0] w_sys_tmp4355;
	wire signed [31:0] w_sys_tmp4356;
	wire signed [31:0] w_sys_tmp4357;
	wire        [31:0] w_sys_tmp4358;
	wire signed [31:0] w_sys_tmp4359;
	wire signed [31:0] w_sys_tmp4360;
	wire signed [31:0] w_sys_tmp4361;
	wire signed [31:0] w_sys_tmp4365;
	wire signed [31:0] w_sys_tmp4368;
	wire        [31:0] w_sys_tmp4369;
	wire signed [31:0] w_sys_tmp4375;
	wire signed [31:0] w_sys_tmp4378;
	wire signed [31:0] w_sys_tmp4379;
	wire signed [31:0] w_sys_tmp4385;
	wire signed [31:0] w_sys_tmp4388;
	wire signed [31:0] w_sys_tmp4395;
	wire signed [31:0] w_sys_tmp4398;
	wire signed [31:0] w_sys_tmp4399;
	wire signed [31:0] w_sys_tmp4405;
	wire signed [31:0] w_sys_tmp4408;
	wire        [31:0] w_sys_tmp4409;
	wire signed [31:0] w_sys_tmp4414;
	wire signed [31:0] w_sys_tmp4793;
	wire               w_sys_tmp4794;
	wire               w_sys_tmp4795;
	wire signed [31:0] w_sys_tmp4796;
	wire signed [31:0] w_sys_tmp4798;
	wire signed [31:0] w_sys_tmp4799;
	wire signed [31:0] w_sys_tmp4801;
	wire signed [31:0] w_sys_tmp4802;
	wire signed [31:0] w_sys_tmp4803;
	wire signed [31:0] w_sys_tmp4804;
	wire        [31:0] w_sys_tmp4805;
	wire signed [31:0] w_sys_tmp4806;
	wire signed [31:0] w_sys_tmp4807;
	wire signed [31:0] w_sys_tmp4808;
	wire signed [31:0] w_sys_tmp4812;
	wire signed [31:0] w_sys_tmp4815;
	wire        [31:0] w_sys_tmp4816;
	wire signed [31:0] w_sys_tmp4822;
	wire signed [31:0] w_sys_tmp4825;
	wire signed [31:0] w_sys_tmp4826;
	wire signed [31:0] w_sys_tmp4832;
	wire signed [31:0] w_sys_tmp4835;
	wire signed [31:0] w_sys_tmp4842;
	wire signed [31:0] w_sys_tmp4845;
	wire signed [31:0] w_sys_tmp4846;
	wire signed [31:0] w_sys_tmp4852;
	wire signed [31:0] w_sys_tmp4855;
	wire        [31:0] w_sys_tmp4856;
	wire signed [31:0] w_sys_tmp4861;
	wire signed [31:0] w_sys_tmp5240;
	wire               w_sys_tmp5241;
	wire               w_sys_tmp5242;
	wire signed [31:0] w_sys_tmp5243;
	wire signed [31:0] w_sys_tmp5245;
	wire signed [31:0] w_sys_tmp5246;
	wire signed [31:0] w_sys_tmp5248;
	wire signed [31:0] w_sys_tmp5249;
	wire signed [31:0] w_sys_tmp5250;
	wire signed [31:0] w_sys_tmp5251;
	wire        [31:0] w_sys_tmp5252;
	wire signed [31:0] w_sys_tmp5253;
	wire signed [31:0] w_sys_tmp5254;
	wire signed [31:0] w_sys_tmp5255;
	wire signed [31:0] w_sys_tmp5259;
	wire signed [31:0] w_sys_tmp5262;
	wire        [31:0] w_sys_tmp5263;
	wire signed [31:0] w_sys_tmp5269;
	wire signed [31:0] w_sys_tmp5272;
	wire signed [31:0] w_sys_tmp5273;
	wire signed [31:0] w_sys_tmp5279;
	wire signed [31:0] w_sys_tmp5282;
	wire signed [31:0] w_sys_tmp5289;
	wire signed [31:0] w_sys_tmp5292;
	wire signed [31:0] w_sys_tmp5293;
	wire signed [31:0] w_sys_tmp5299;
	wire signed [31:0] w_sys_tmp5302;
	wire        [31:0] w_sys_tmp5303;
	wire signed [31:0] w_sys_tmp5308;
	wire signed [31:0] w_sys_tmp5687;
	wire               w_sys_tmp5688;
	wire               w_sys_tmp5689;
	wire signed [31:0] w_sys_tmp5690;
	wire signed [31:0] w_sys_tmp5691;
	wire signed [31:0] w_sys_tmp5692;
	wire               w_sys_tmp5693;
	wire               w_sys_tmp5694;
	wire signed [31:0] w_sys_tmp5695;
	wire signed [31:0] w_sys_tmp5698;
	wire signed [31:0] w_sys_tmp5699;
	wire signed [31:0] w_sys_tmp5700;
	wire        [31:0] w_sys_tmp5701;
	wire signed [31:0] w_sys_tmp5702;
	wire signed [31:0] w_sys_tmp5703;
	wire signed [31:0] w_sys_tmp5705;
	wire signed [31:0] w_sys_tmp5706;
	wire signed [31:0] w_sys_tmp5767;
	wire               w_sys_tmp5768;
	wire               w_sys_tmp5769;
	wire signed [31:0] w_sys_tmp5770;
	wire signed [31:0] w_sys_tmp5772;
	wire signed [31:0] w_sys_tmp5773;
	wire signed [31:0] w_sys_tmp5775;
	wire signed [31:0] w_sys_tmp5776;
	wire signed [31:0] w_sys_tmp5777;
	wire        [31:0] w_sys_tmp5778;
	wire signed [31:0] w_sys_tmp5779;
	wire signed [31:0] w_sys_tmp5780;
	wire signed [31:0] w_sys_tmp5782;
	wire signed [31:0] w_sys_tmp5783;
	wire signed [31:0] w_sys_tmp5784;
	wire signed [31:0] w_sys_tmp5863;
	wire               w_sys_tmp5864;
	wire               w_sys_tmp5865;
	wire signed [31:0] w_sys_tmp5866;
	wire signed [31:0] w_sys_tmp5868;
	wire signed [31:0] w_sys_tmp5869;
	wire signed [31:0] w_sys_tmp5871;
	wire signed [31:0] w_sys_tmp5872;
	wire signed [31:0] w_sys_tmp5873;
	wire        [31:0] w_sys_tmp5874;
	wire signed [31:0] w_sys_tmp5875;
	wire signed [31:0] w_sys_tmp5876;
	wire signed [31:0] w_sys_tmp5878;
	wire signed [31:0] w_sys_tmp5879;
	wire signed [31:0] w_sys_tmp5880;
	wire signed [31:0] w_sys_tmp5959;
	wire               w_sys_tmp5960;
	wire               w_sys_tmp5961;
	wire signed [31:0] w_sys_tmp5962;
	wire signed [31:0] w_sys_tmp5964;
	wire signed [31:0] w_sys_tmp5965;
	wire signed [31:0] w_sys_tmp5967;
	wire signed [31:0] w_sys_tmp5968;
	wire signed [31:0] w_sys_tmp5969;
	wire        [31:0] w_sys_tmp5970;
	wire signed [31:0] w_sys_tmp5971;
	wire signed [31:0] w_sys_tmp5972;
	wire signed [31:0] w_sys_tmp5974;
	wire signed [31:0] w_sys_tmp5975;
	wire signed [31:0] w_sys_tmp5976;
	wire signed [31:0] w_sys_tmp6055;
	wire               w_sys_tmp6056;
	wire               w_sys_tmp6057;
	wire signed [31:0] w_sys_tmp6058;
	wire signed [31:0] w_sys_tmp6059;
	wire signed [31:0] w_sys_tmp6060;
	wire               w_sys_tmp6061;
	wire               w_sys_tmp6062;
	wire signed [31:0] w_sys_tmp6063;
	wire signed [31:0] w_sys_tmp6066;
	wire signed [31:0] w_sys_tmp6067;
	wire signed [31:0] w_sys_tmp6068;
	wire        [31:0] w_sys_tmp6069;
	wire signed [31:0] w_sys_tmp6070;
	wire signed [31:0] w_sys_tmp6071;
	wire signed [31:0] w_sys_tmp6073;
	wire signed [31:0] w_sys_tmp6074;
	wire signed [31:0] w_sys_tmp6135;
	wire               w_sys_tmp6136;
	wire               w_sys_tmp6137;
	wire signed [31:0] w_sys_tmp6138;
	wire signed [31:0] w_sys_tmp6140;
	wire signed [31:0] w_sys_tmp6141;
	wire signed [31:0] w_sys_tmp6143;
	wire signed [31:0] w_sys_tmp6144;
	wire signed [31:0] w_sys_tmp6145;
	wire        [31:0] w_sys_tmp6146;
	wire signed [31:0] w_sys_tmp6147;
	wire signed [31:0] w_sys_tmp6148;
	wire signed [31:0] w_sys_tmp6150;
	wire signed [31:0] w_sys_tmp6151;
	wire signed [31:0] w_sys_tmp6152;
	wire signed [31:0] w_sys_tmp6231;
	wire               w_sys_tmp6232;
	wire               w_sys_tmp6233;
	wire signed [31:0] w_sys_tmp6234;
	wire signed [31:0] w_sys_tmp6236;
	wire signed [31:0] w_sys_tmp6237;
	wire signed [31:0] w_sys_tmp6239;
	wire signed [31:0] w_sys_tmp6240;
	wire signed [31:0] w_sys_tmp6241;
	wire        [31:0] w_sys_tmp6242;
	wire signed [31:0] w_sys_tmp6243;
	wire signed [31:0] w_sys_tmp6244;
	wire signed [31:0] w_sys_tmp6246;
	wire signed [31:0] w_sys_tmp6247;
	wire signed [31:0] w_sys_tmp6248;
	wire signed [31:0] w_sys_tmp6327;
	wire               w_sys_tmp6328;
	wire               w_sys_tmp6329;
	wire signed [31:0] w_sys_tmp6330;
	wire signed [31:0] w_sys_tmp6332;
	wire signed [31:0] w_sys_tmp6333;
	wire signed [31:0] w_sys_tmp6335;
	wire signed [31:0] w_sys_tmp6336;
	wire signed [31:0] w_sys_tmp6337;
	wire        [31:0] w_sys_tmp6338;
	wire signed [31:0] w_sys_tmp6339;
	wire signed [31:0] w_sys_tmp6340;
	wire signed [31:0] w_sys_tmp6342;
	wire signed [31:0] w_sys_tmp6343;
	wire signed [31:0] w_sys_tmp6344;
	wire signed [31:0] w_sys_tmp6423;
	wire               w_sys_tmp6424;
	wire               w_sys_tmp6425;
	wire signed [31:0] w_sys_tmp6426;
	wire signed [31:0] w_sys_tmp6427;
	wire signed [31:0] w_sys_tmp6428;
	wire               w_sys_tmp6429;
	wire               w_sys_tmp6430;
	wire signed [31:0] w_sys_tmp6431;
	wire signed [31:0] w_sys_tmp6434;
	wire signed [31:0] w_sys_tmp6435;
	wire signed [31:0] w_sys_tmp6436;
	wire        [31:0] w_sys_tmp6437;
	wire signed [31:0] w_sys_tmp6438;
	wire signed [31:0] w_sys_tmp6439;
	wire signed [31:0] w_sys_tmp6441;
	wire signed [31:0] w_sys_tmp6442;
	wire signed [31:0] w_sys_tmp6503;
	wire               w_sys_tmp6504;
	wire               w_sys_tmp6505;
	wire signed [31:0] w_sys_tmp6506;
	wire signed [31:0] w_sys_tmp6508;
	wire signed [31:0] w_sys_tmp6509;
	wire signed [31:0] w_sys_tmp6511;
	wire signed [31:0] w_sys_tmp6512;
	wire signed [31:0] w_sys_tmp6513;
	wire        [31:0] w_sys_tmp6514;
	wire signed [31:0] w_sys_tmp6515;
	wire signed [31:0] w_sys_tmp6516;
	wire signed [31:0] w_sys_tmp6518;
	wire signed [31:0] w_sys_tmp6519;
	wire signed [31:0] w_sys_tmp6520;
	wire signed [31:0] w_sys_tmp6599;
	wire               w_sys_tmp6600;
	wire               w_sys_tmp6601;
	wire signed [31:0] w_sys_tmp6602;
	wire signed [31:0] w_sys_tmp6604;
	wire signed [31:0] w_sys_tmp6605;
	wire signed [31:0] w_sys_tmp6607;
	wire signed [31:0] w_sys_tmp6608;
	wire signed [31:0] w_sys_tmp6609;
	wire        [31:0] w_sys_tmp6610;
	wire signed [31:0] w_sys_tmp6611;
	wire signed [31:0] w_sys_tmp6612;
	wire signed [31:0] w_sys_tmp6614;
	wire signed [31:0] w_sys_tmp6615;
	wire signed [31:0] w_sys_tmp6616;
	wire signed [31:0] w_sys_tmp6695;
	wire               w_sys_tmp6696;
	wire               w_sys_tmp6697;
	wire signed [31:0] w_sys_tmp6698;
	wire signed [31:0] w_sys_tmp6700;
	wire signed [31:0] w_sys_tmp6701;
	wire signed [31:0] w_sys_tmp6703;
	wire signed [31:0] w_sys_tmp6704;
	wire signed [31:0] w_sys_tmp6705;
	wire        [31:0] w_sys_tmp6706;
	wire signed [31:0] w_sys_tmp6707;
	wire signed [31:0] w_sys_tmp6708;
	wire signed [31:0] w_sys_tmp6710;
	wire signed [31:0] w_sys_tmp6711;
	wire signed [31:0] w_sys_tmp6712;
	wire signed [31:0] w_sys_tmp6791;
	wire               w_sys_tmp6792;
	wire               w_sys_tmp6793;
	wire signed [31:0] w_sys_tmp6794;
	wire signed [31:0] w_sys_tmp6795;
	wire signed [31:0] w_sys_tmp6796;
	wire               w_sys_tmp6797;
	wire               w_sys_tmp6798;
	wire signed [31:0] w_sys_tmp6799;
	wire signed [31:0] w_sys_tmp6802;
	wire signed [31:0] w_sys_tmp6803;
	wire signed [31:0] w_sys_tmp6804;
	wire        [31:0] w_sys_tmp6805;
	wire signed [31:0] w_sys_tmp6806;
	wire signed [31:0] w_sys_tmp6807;
	wire signed [31:0] w_sys_tmp6809;
	wire signed [31:0] w_sys_tmp6810;
	wire signed [31:0] w_sys_tmp6871;
	wire               w_sys_tmp6872;
	wire               w_sys_tmp6873;
	wire signed [31:0] w_sys_tmp6874;
	wire signed [31:0] w_sys_tmp6876;
	wire signed [31:0] w_sys_tmp6877;
	wire signed [31:0] w_sys_tmp6879;
	wire signed [31:0] w_sys_tmp6880;
	wire signed [31:0] w_sys_tmp6881;
	wire        [31:0] w_sys_tmp6882;
	wire signed [31:0] w_sys_tmp6883;
	wire signed [31:0] w_sys_tmp6884;
	wire signed [31:0] w_sys_tmp6886;
	wire signed [31:0] w_sys_tmp6887;
	wire signed [31:0] w_sys_tmp6888;
	wire signed [31:0] w_sys_tmp6967;
	wire               w_sys_tmp6968;
	wire               w_sys_tmp6969;
	wire signed [31:0] w_sys_tmp6970;
	wire signed [31:0] w_sys_tmp6972;
	wire signed [31:0] w_sys_tmp6973;
	wire signed [31:0] w_sys_tmp6975;
	wire signed [31:0] w_sys_tmp6976;
	wire signed [31:0] w_sys_tmp6977;
	wire        [31:0] w_sys_tmp6978;
	wire signed [31:0] w_sys_tmp6979;
	wire signed [31:0] w_sys_tmp6980;
	wire signed [31:0] w_sys_tmp6982;
	wire signed [31:0] w_sys_tmp6983;
	wire signed [31:0] w_sys_tmp6984;
	wire signed [31:0] w_sys_tmp7063;
	wire               w_sys_tmp7064;
	wire               w_sys_tmp7065;
	wire signed [31:0] w_sys_tmp7066;
	wire signed [31:0] w_sys_tmp7068;
	wire signed [31:0] w_sys_tmp7069;
	wire signed [31:0] w_sys_tmp7071;
	wire signed [31:0] w_sys_tmp7072;
	wire signed [31:0] w_sys_tmp7073;
	wire        [31:0] w_sys_tmp7074;
	wire signed [31:0] w_sys_tmp7075;
	wire signed [31:0] w_sys_tmp7076;
	wire signed [31:0] w_sys_tmp7078;
	wire signed [31:0] w_sys_tmp7079;
	wire signed [31:0] w_sys_tmp7080;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign w_fld_T_0_addr_0 = 15'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 15'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 15'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_fld_V_3_addr_0 = 15'sh0;
	assign w_fld_V_3_datain_0 = 32'h0;
	assign w_fld_V_3_r_w_0 = 1'h0;
	assign w_fld_V_3_ce_0 = w_sys_ce;
	assign w_fld_V_3_ce_1 = w_sys_ce;
	assign w_sub09_T_addr = ( (|r_sys_processing_methodID) ? r_sub09_T_addr : 15'sh0 ) ;
	assign w_sub09_T_datain = ( (|r_sys_processing_methodID) ? r_sub09_T_datain : 32'h0 ) ;
	assign w_sub09_T_r_w = ( (|r_sys_processing_methodID) ? r_sub09_T_r_w : 1'h0 ) ;
	assign w_sub09_V_addr = ( (|r_sys_processing_methodID) ? r_sub09_V_addr : 15'sh0 ) ;
	assign w_sub09_V_datain = ( (|r_sys_processing_methodID) ? r_sub09_V_datain : 32'h0 ) ;
	assign w_sub09_V_r_w = ( (|r_sys_processing_methodID) ? r_sub09_V_r_w : 1'h0 ) ;
	assign w_sub09_U_addr = ( (|r_sys_processing_methodID) ? r_sub09_U_addr : 15'sh0 ) ;
	assign w_sub09_U_datain = ( (|r_sys_processing_methodID) ? r_sub09_U_datain : 32'h0 ) ;
	assign w_sub09_U_r_w = ( (|r_sys_processing_methodID) ? r_sub09_U_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 15'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_T_addr = ( (|r_sys_processing_methodID) ? r_sub08_T_addr : 15'sh0 ) ;
	assign w_sub08_T_datain = ( (|r_sys_processing_methodID) ? r_sub08_T_datain : 32'h0 ) ;
	assign w_sub08_T_r_w = ( (|r_sys_processing_methodID) ? r_sub08_T_r_w : 1'h0 ) ;
	assign w_sub08_V_addr = ( (|r_sys_processing_methodID) ? r_sub08_V_addr : 15'sh0 ) ;
	assign w_sub08_V_datain = ( (|r_sys_processing_methodID) ? r_sub08_V_datain : 32'h0 ) ;
	assign w_sub08_V_r_w = ( (|r_sys_processing_methodID) ? r_sub08_V_r_w : 1'h0 ) ;
	assign w_sub08_U_addr = ( (|r_sys_processing_methodID) ? r_sub08_U_addr : 15'sh0 ) ;
	assign w_sub08_U_datain = ( (|r_sys_processing_methodID) ? r_sub08_U_datain : 32'h0 ) ;
	assign w_sub08_U_r_w = ( (|r_sys_processing_methodID) ? r_sub08_U_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 15'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub12_T_addr = ( (|r_sys_processing_methodID) ? r_sub12_T_addr : 15'sh0 ) ;
	assign w_sub12_T_datain = ( (|r_sys_processing_methodID) ? r_sub12_T_datain : 32'h0 ) ;
	assign w_sub12_T_r_w = ( (|r_sys_processing_methodID) ? r_sub12_T_r_w : 1'h0 ) ;
	assign w_sub12_V_addr = ( (|r_sys_processing_methodID) ? r_sub12_V_addr : 15'sh0 ) ;
	assign w_sub12_V_datain = ( (|r_sys_processing_methodID) ? r_sub12_V_datain : 32'h0 ) ;
	assign w_sub12_V_r_w = ( (|r_sys_processing_methodID) ? r_sub12_V_r_w : 1'h0 ) ;
	assign w_sub12_U_addr = ( (|r_sys_processing_methodID) ? r_sub12_U_addr : 15'sh0 ) ;
	assign w_sub12_U_datain = ( (|r_sys_processing_methodID) ? r_sub12_U_datain : 32'h0 ) ;
	assign w_sub12_U_r_w = ( (|r_sys_processing_methodID) ? r_sub12_U_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 15'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_T_addr = ( (|r_sys_processing_methodID) ? r_sub03_T_addr : 15'sh0 ) ;
	assign w_sub03_T_datain = ( (|r_sys_processing_methodID) ? r_sub03_T_datain : 32'h0 ) ;
	assign w_sub03_T_r_w = ( (|r_sys_processing_methodID) ? r_sub03_T_r_w : 1'h0 ) ;
	assign w_sub03_V_addr = ( (|r_sys_processing_methodID) ? r_sub03_V_addr : 15'sh0 ) ;
	assign w_sub03_V_datain = ( (|r_sys_processing_methodID) ? r_sub03_V_datain : 32'h0 ) ;
	assign w_sub03_V_r_w = ( (|r_sys_processing_methodID) ? r_sub03_V_r_w : 1'h0 ) ;
	assign w_sub03_U_addr = ( (|r_sys_processing_methodID) ? r_sub03_U_addr : 15'sh0 ) ;
	assign w_sub03_U_datain = ( (|r_sys_processing_methodID) ? r_sub03_U_datain : 32'h0 ) ;
	assign w_sub03_U_r_w = ( (|r_sys_processing_methodID) ? r_sub03_U_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 15'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_T_addr = ( (|r_sys_processing_methodID) ? r_sub02_T_addr : 15'sh0 ) ;
	assign w_sub02_T_datain = ( (|r_sys_processing_methodID) ? r_sub02_T_datain : 32'h0 ) ;
	assign w_sub02_T_r_w = ( (|r_sys_processing_methodID) ? r_sub02_T_r_w : 1'h0 ) ;
	assign w_sub02_V_addr = ( (|r_sys_processing_methodID) ? r_sub02_V_addr : 15'sh0 ) ;
	assign w_sub02_V_datain = ( (|r_sys_processing_methodID) ? r_sub02_V_datain : 32'h0 ) ;
	assign w_sub02_V_r_w = ( (|r_sys_processing_methodID) ? r_sub02_V_r_w : 1'h0 ) ;
	assign w_sub02_U_addr = ( (|r_sys_processing_methodID) ? r_sub02_U_addr : 15'sh0 ) ;
	assign w_sub02_U_datain = ( (|r_sys_processing_methodID) ? r_sub02_U_datain : 32'h0 ) ;
	assign w_sub02_U_r_w = ( (|r_sys_processing_methodID) ? r_sub02_U_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 15'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_T_addr = ( (|r_sys_processing_methodID) ? r_sub11_T_addr : 15'sh0 ) ;
	assign w_sub11_T_datain = ( (|r_sys_processing_methodID) ? r_sub11_T_datain : 32'h0 ) ;
	assign w_sub11_T_r_w = ( (|r_sys_processing_methodID) ? r_sub11_T_r_w : 1'h0 ) ;
	assign w_sub11_V_addr = ( (|r_sys_processing_methodID) ? r_sub11_V_addr : 15'sh0 ) ;
	assign w_sub11_V_datain = ( (|r_sys_processing_methodID) ? r_sub11_V_datain : 32'h0 ) ;
	assign w_sub11_V_r_w = ( (|r_sys_processing_methodID) ? r_sub11_V_r_w : 1'h0 ) ;
	assign w_sub11_U_addr = ( (|r_sys_processing_methodID) ? r_sub11_U_addr : 15'sh0 ) ;
	assign w_sub11_U_datain = ( (|r_sys_processing_methodID) ? r_sub11_U_datain : 32'h0 ) ;
	assign w_sub11_U_r_w = ( (|r_sys_processing_methodID) ? r_sub11_U_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 15'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_T_addr = ( (|r_sys_processing_methodID) ? r_sub14_T_addr : 15'sh0 ) ;
	assign w_sub14_T_datain = ( (|r_sys_processing_methodID) ? r_sub14_T_datain : 32'h0 ) ;
	assign w_sub14_T_r_w = ( (|r_sys_processing_methodID) ? r_sub14_T_r_w : 1'h0 ) ;
	assign w_sub14_V_addr = ( (|r_sys_processing_methodID) ? r_sub14_V_addr : 15'sh0 ) ;
	assign w_sub14_V_datain = ( (|r_sys_processing_methodID) ? r_sub14_V_datain : 32'h0 ) ;
	assign w_sub14_V_r_w = ( (|r_sys_processing_methodID) ? r_sub14_V_r_w : 1'h0 ) ;
	assign w_sub14_U_addr = ( (|r_sys_processing_methodID) ? r_sub14_U_addr : 15'sh0 ) ;
	assign w_sub14_U_datain = ( (|r_sys_processing_methodID) ? r_sub14_U_datain : 32'h0 ) ;
	assign w_sub14_U_r_w = ( (|r_sys_processing_methodID) ? r_sub14_U_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 15'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_T_addr = ( (|r_sys_processing_methodID) ? r_sub01_T_addr : 15'sh0 ) ;
	assign w_sub01_T_datain = ( (|r_sys_processing_methodID) ? r_sub01_T_datain : 32'h0 ) ;
	assign w_sub01_T_r_w = ( (|r_sys_processing_methodID) ? r_sub01_T_r_w : 1'h0 ) ;
	assign w_sub01_V_addr = ( (|r_sys_processing_methodID) ? r_sub01_V_addr : 15'sh0 ) ;
	assign w_sub01_V_datain = ( (|r_sys_processing_methodID) ? r_sub01_V_datain : 32'h0 ) ;
	assign w_sub01_V_r_w = ( (|r_sys_processing_methodID) ? r_sub01_V_r_w : 1'h0 ) ;
	assign w_sub01_U_addr = ( (|r_sys_processing_methodID) ? r_sub01_U_addr : 15'sh0 ) ;
	assign w_sub01_U_datain = ( (|r_sys_processing_methodID) ? r_sub01_U_datain : 32'h0 ) ;
	assign w_sub01_U_r_w = ( (|r_sys_processing_methodID) ? r_sub01_U_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 15'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub13_T_addr = ( (|r_sys_processing_methodID) ? r_sub13_T_addr : 15'sh0 ) ;
	assign w_sub13_T_datain = ( (|r_sys_processing_methodID) ? r_sub13_T_datain : 32'h0 ) ;
	assign w_sub13_T_r_w = ( (|r_sys_processing_methodID) ? r_sub13_T_r_w : 1'h0 ) ;
	assign w_sub13_V_addr = ( (|r_sys_processing_methodID) ? r_sub13_V_addr : 15'sh0 ) ;
	assign w_sub13_V_datain = ( (|r_sys_processing_methodID) ? r_sub13_V_datain : 32'h0 ) ;
	assign w_sub13_V_r_w = ( (|r_sys_processing_methodID) ? r_sub13_V_r_w : 1'h0 ) ;
	assign w_sub13_U_addr = ( (|r_sys_processing_methodID) ? r_sub13_U_addr : 15'sh0 ) ;
	assign w_sub13_U_datain = ( (|r_sys_processing_methodID) ? r_sub13_U_datain : 32'h0 ) ;
	assign w_sub13_U_r_w = ( (|r_sys_processing_methodID) ? r_sub13_U_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 15'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub00_T_addr = ( (|r_sys_processing_methodID) ? r_sub00_T_addr : 15'sh0 ) ;
	assign w_sub00_T_datain = ( (|r_sys_processing_methodID) ? r_sub00_T_datain : 32'h0 ) ;
	assign w_sub00_T_r_w = ( (|r_sys_processing_methodID) ? r_sub00_T_r_w : 1'h0 ) ;
	assign w_sub00_V_addr = ( (|r_sys_processing_methodID) ? r_sub00_V_addr : 15'sh0 ) ;
	assign w_sub00_V_datain = ( (|r_sys_processing_methodID) ? r_sub00_V_datain : 32'h0 ) ;
	assign w_sub00_V_r_w = ( (|r_sys_processing_methodID) ? r_sub00_V_r_w : 1'h0 ) ;
	assign w_sub00_U_addr = ( (|r_sys_processing_methodID) ? r_sub00_U_addr : 15'sh0 ) ;
	assign w_sub00_U_datain = ( (|r_sys_processing_methodID) ? r_sub00_U_datain : 32'h0 ) ;
	assign w_sub00_U_r_w = ( (|r_sys_processing_methodID) ? r_sub00_U_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 15'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_T_addr = ( (|r_sys_processing_methodID) ? r_sub07_T_addr : 15'sh0 ) ;
	assign w_sub07_T_datain = ( (|r_sys_processing_methodID) ? r_sub07_T_datain : 32'h0 ) ;
	assign w_sub07_T_r_w = ( (|r_sys_processing_methodID) ? r_sub07_T_r_w : 1'h0 ) ;
	assign w_sub07_V_addr = ( (|r_sys_processing_methodID) ? r_sub07_V_addr : 15'sh0 ) ;
	assign w_sub07_V_datain = ( (|r_sys_processing_methodID) ? r_sub07_V_datain : 32'h0 ) ;
	assign w_sub07_V_r_w = ( (|r_sys_processing_methodID) ? r_sub07_V_r_w : 1'h0 ) ;
	assign w_sub07_U_addr = ( (|r_sys_processing_methodID) ? r_sub07_U_addr : 15'sh0 ) ;
	assign w_sub07_U_datain = ( (|r_sys_processing_methodID) ? r_sub07_U_datain : 32'h0 ) ;
	assign w_sub07_U_r_w = ( (|r_sys_processing_methodID) ? r_sub07_U_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 15'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_T_addr = ( (|r_sys_processing_methodID) ? r_sub06_T_addr : 15'sh0 ) ;
	assign w_sub06_T_datain = ( (|r_sys_processing_methodID) ? r_sub06_T_datain : 32'h0 ) ;
	assign w_sub06_T_r_w = ( (|r_sys_processing_methodID) ? r_sub06_T_r_w : 1'h0 ) ;
	assign w_sub06_V_addr = ( (|r_sys_processing_methodID) ? r_sub06_V_addr : 15'sh0 ) ;
	assign w_sub06_V_datain = ( (|r_sys_processing_methodID) ? r_sub06_V_datain : 32'h0 ) ;
	assign w_sub06_V_r_w = ( (|r_sys_processing_methodID) ? r_sub06_V_r_w : 1'h0 ) ;
	assign w_sub06_U_addr = ( (|r_sys_processing_methodID) ? r_sub06_U_addr : 15'sh0 ) ;
	assign w_sub06_U_datain = ( (|r_sys_processing_methodID) ? r_sub06_U_datain : 32'h0 ) ;
	assign w_sub06_U_r_w = ( (|r_sys_processing_methodID) ? r_sub06_U_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 15'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_T_addr = ( (|r_sys_processing_methodID) ? r_sub15_T_addr : 15'sh0 ) ;
	assign w_sub15_T_datain = ( (|r_sys_processing_methodID) ? r_sub15_T_datain : 32'h0 ) ;
	assign w_sub15_T_r_w = ( (|r_sys_processing_methodID) ? r_sub15_T_r_w : 1'h0 ) ;
	assign w_sub15_V_addr = ( (|r_sys_processing_methodID) ? r_sub15_V_addr : 15'sh0 ) ;
	assign w_sub15_V_datain = ( (|r_sys_processing_methodID) ? r_sub15_V_datain : 32'h0 ) ;
	assign w_sub15_V_r_w = ( (|r_sys_processing_methodID) ? r_sub15_V_r_w : 1'h0 ) ;
	assign w_sub15_U_addr = ( (|r_sys_processing_methodID) ? r_sub15_U_addr : 15'sh0 ) ;
	assign w_sub15_U_datain = ( (|r_sys_processing_methodID) ? r_sub15_U_datain : 32'h0 ) ;
	assign w_sub15_U_r_w = ( (|r_sys_processing_methodID) ? r_sub15_U_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 15'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_T_addr = ( (|r_sys_processing_methodID) ? r_sub05_T_addr : 15'sh0 ) ;
	assign w_sub05_T_datain = ( (|r_sys_processing_methodID) ? r_sub05_T_datain : 32'h0 ) ;
	assign w_sub05_T_r_w = ( (|r_sys_processing_methodID) ? r_sub05_T_r_w : 1'h0 ) ;
	assign w_sub05_V_addr = ( (|r_sys_processing_methodID) ? r_sub05_V_addr : 15'sh0 ) ;
	assign w_sub05_V_datain = ( (|r_sys_processing_methodID) ? r_sub05_V_datain : 32'h0 ) ;
	assign w_sub05_V_r_w = ( (|r_sys_processing_methodID) ? r_sub05_V_r_w : 1'h0 ) ;
	assign w_sub05_U_addr = ( (|r_sys_processing_methodID) ? r_sub05_U_addr : 15'sh0 ) ;
	assign w_sub05_U_datain = ( (|r_sys_processing_methodID) ? r_sub05_U_datain : 32'h0 ) ;
	assign w_sub05_U_r_w = ( (|r_sys_processing_methodID) ? r_sub05_U_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 15'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_T_addr = ( (|r_sys_processing_methodID) ? r_sub04_T_addr : 15'sh0 ) ;
	assign w_sub04_T_datain = ( (|r_sys_processing_methodID) ? r_sub04_T_datain : 32'h0 ) ;
	assign w_sub04_T_r_w = ( (|r_sys_processing_methodID) ? r_sub04_T_r_w : 1'h0 ) ;
	assign w_sub04_V_addr = ( (|r_sys_processing_methodID) ? r_sub04_V_addr : 15'sh0 ) ;
	assign w_sub04_V_datain = ( (|r_sys_processing_methodID) ? r_sub04_V_datain : 32'h0 ) ;
	assign w_sub04_V_r_w = ( (|r_sys_processing_methodID) ? r_sub04_V_r_w : 1'h0 ) ;
	assign w_sub04_U_addr = ( (|r_sys_processing_methodID) ? r_sub04_U_addr : 15'sh0 ) ;
	assign w_sub04_U_datain = ( (|r_sys_processing_methodID) ? r_sub04_U_datain : 32'h0 ) ;
	assign w_sub04_U_r_w = ( (|r_sys_processing_methodID) ? r_sub04_U_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 15'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_T_addr = ( (|r_sys_processing_methodID) ? r_sub10_T_addr : 15'sh0 ) ;
	assign w_sub10_T_datain = ( (|r_sys_processing_methodID) ? r_sub10_T_datain : 32'h0 ) ;
	assign w_sub10_T_r_w = ( (|r_sys_processing_methodID) ? r_sub10_T_r_w : 1'h0 ) ;
	assign w_sub10_V_addr = ( (|r_sys_processing_methodID) ? r_sub10_V_addr : 15'sh0 ) ;
	assign w_sub10_V_datain = ( (|r_sys_processing_methodID) ? r_sub10_V_datain : 32'h0 ) ;
	assign w_sub10_V_r_w = ( (|r_sys_processing_methodID) ? r_sub10_V_r_w : 1'h0 ) ;
	assign w_sub10_U_addr = ( (|r_sys_processing_methodID) ? r_sub10_U_addr : 15'sh0 ) ;
	assign w_sub10_U_datain = ( (|r_sys_processing_methodID) ? r_sub10_U_datain : 32'h0 ) ;
	assign w_sub10_U_r_w = ( (|r_sys_processing_methodID) ? r_sub10_U_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 15'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000080;
	assign w_sys_tmp3 = 32'sh00000081;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'sh00000002;
	assign w_sys_tmp7 = 32'h3d000000;
	assign w_sys_tmp8 = 32'h3c000000;
	assign w_sys_tmp9 = 32'h3c03126f;
	assign w_sys_tmp10 = 32'h3d03126f;
	assign w_sys_tmp11 = 32'h3f03126f;
	assign w_sys_tmp12 = 32'h4103126f;
	assign w_sys_tmp13 = ( !w_sys_tmp14 );
	assign w_sys_tmp14 = (r_run_my_24 < r_run_k_20);
	assign w_sys_tmp15 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp16 = ( !w_sys_tmp17 );
	assign w_sys_tmp17 = (r_run_mx_23 < r_run_j_21);
	assign w_sys_tmp19 = w_ip_MultFloat_product_0;
	assign w_sys_tmp20 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp21 = (r_run_k_20 - w_sys_intOne);
	assign w_sys_tmp23 = (w_sys_tmp24 + r_run_k_20);
	assign w_sys_tmp24 = (r_run_j_21 * w_sys_tmp25);
	assign w_sys_tmp25 = 32'sh00000081;
	assign w_sys_tmp26 = 32'h0;
	assign w_sys_tmp28 = (w_sys_tmp29 + r_run_k_20);
	assign w_sys_tmp29 = (r_run_copy2_j_39 * w_sys_tmp25);
	assign w_sys_tmp33 = (w_sys_tmp34 + r_run_k_20);
	assign w_sys_tmp34 = (r_run_copy1_j_38 * w_sys_tmp25);
	assign w_sys_tmp37 = 32'h42200000;
	assign w_sys_tmp38 = w_sys_tmp19;
	assign w_sys_tmp39 = 32'h3f800000;
	assign w_sys_tmp42 = (w_sys_tmp43 + r_run_k_20);
	assign w_sys_tmp43 = (r_run_copy0_j_37 * w_sys_tmp25);
	assign w_sys_tmp46 = (r_run_copy0_j_37 + w_sys_intOne);
	assign w_sys_tmp47 = (r_run_copy1_j_38 + w_sys_intOne);
	assign w_sys_tmp48 = (r_run_copy2_j_39 + w_sys_intOne);
	assign w_sys_tmp49 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp129 = r_sys_tmp4_float;
	assign w_sys_tmp227 = ( !w_sys_tmp228 );
	assign w_sys_tmp228 = (w_sys_tmp229 < r_run_k_20);
	assign w_sys_tmp229 = 32'sh00000021;
	assign w_sys_tmp230 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp231 = ( !w_sys_tmp232 );
	assign w_sys_tmp232 = (w_sys_tmp233 < r_run_j_21);
	assign w_sys_tmp233 = 32'sh00000021;
	assign w_sys_tmp236 = (w_sys_tmp237 + r_run_k_20);
	assign w_sys_tmp237 = (r_run_j_21 * w_sys_tmp238);
	assign w_sys_tmp238 = 32'sh00000081;
	assign w_sys_tmp239 = w_fld_U_2_dataout_1;
	assign w_sys_tmp240 = (w_sys_tmp241 + r_run_k_20);
	assign w_sys_tmp241 = (r_run_copy4_j_44 * w_sys_tmp238);
	assign w_sys_tmp244 = (w_sys_tmp245 + r_run_k_20);
	assign w_sys_tmp245 = (r_run_copy3_j_43 * w_sys_tmp238);
	assign w_sys_tmp247 = w_fld_V_3_dataout_1;
	assign w_sys_tmp248 = (w_sys_tmp249 + r_run_k_20);
	assign w_sys_tmp249 = (r_run_copy2_j_42 * w_sys_tmp238);
	assign w_sys_tmp252 = (w_sys_tmp253 + r_run_k_20);
	assign w_sys_tmp253 = (r_run_copy1_j_41 * w_sys_tmp238);
	assign w_sys_tmp255 = w_fld_T_0_dataout_1;
	assign w_sys_tmp256 = (w_sys_tmp257 + r_run_k_20);
	assign w_sys_tmp257 = (r_run_copy0_j_40 * w_sys_tmp238);
	assign w_sys_tmp259 = (r_run_copy0_j_40 + w_sys_intOne);
	assign w_sys_tmp260 = (r_run_copy1_j_41 + w_sys_intOne);
	assign w_sys_tmp261 = (r_run_copy2_j_42 + w_sys_intOne);
	assign w_sys_tmp262 = (r_run_copy3_j_43 + w_sys_intOne);
	assign w_sys_tmp263 = (r_run_copy4_j_44 + w_sys_intOne);
	assign w_sys_tmp264 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp445 = 32'sh00000020;
	assign w_sys_tmp446 = ( !w_sys_tmp447 );
	assign w_sys_tmp447 = (w_sys_tmp448 < r_run_j_21);
	assign w_sys_tmp448 = 32'sh00000041;
	assign w_sys_tmp451 = (w_sys_tmp452 + r_run_k_20);
	assign w_sys_tmp452 = (r_run_j_21 * w_sys_tmp453);
	assign w_sys_tmp453 = 32'sh00000081;
	assign w_sys_tmp454 = w_fld_U_2_dataout_1;
	assign w_sys_tmp455 = (w_sys_tmp456 + r_run_k_20);
	assign w_sys_tmp456 = (r_run_copy4_j_49 * w_sys_tmp453);
	assign w_sys_tmp459 = (w_sys_tmp460 + r_run_k_20);
	assign w_sys_tmp460 = (r_run_copy3_j_48 * w_sys_tmp453);
	assign w_sys_tmp462 = w_fld_V_3_dataout_1;
	assign w_sys_tmp463 = (w_sys_tmp464 + r_run_k_20);
	assign w_sys_tmp464 = (r_run_copy2_j_47 * w_sys_tmp453);
	assign w_sys_tmp467 = (w_sys_tmp468 + r_run_k_20);
	assign w_sys_tmp468 = (r_run_copy1_j_46 * w_sys_tmp453);
	assign w_sys_tmp470 = w_fld_T_0_dataout_1;
	assign w_sys_tmp471 = (w_sys_tmp472 + r_run_k_20);
	assign w_sys_tmp472 = (r_run_copy0_j_45 * w_sys_tmp453);
	assign w_sys_tmp474 = (r_run_copy0_j_45 + w_sys_intOne);
	assign w_sys_tmp475 = (r_run_copy1_j_46 + w_sys_intOne);
	assign w_sys_tmp476 = (r_run_copy2_j_47 + w_sys_intOne);
	assign w_sys_tmp477 = (r_run_copy3_j_48 + w_sys_intOne);
	assign w_sys_tmp478 = (r_run_copy4_j_49 + w_sys_intOne);
	assign w_sys_tmp479 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp660 = 32'sh00000040;
	assign w_sys_tmp661 = ( !w_sys_tmp662 );
	assign w_sys_tmp662 = (w_sys_tmp663 < r_run_j_21);
	assign w_sys_tmp663 = 32'sh00000061;
	assign w_sys_tmp666 = (w_sys_tmp667 + r_run_k_20);
	assign w_sys_tmp667 = (r_run_j_21 * w_sys_tmp668);
	assign w_sys_tmp668 = 32'sh00000081;
	assign w_sys_tmp669 = w_fld_U_2_dataout_1;
	assign w_sys_tmp670 = (w_sys_tmp671 + r_run_k_20);
	assign w_sys_tmp671 = (r_run_copy4_j_54 * w_sys_tmp668);
	assign w_sys_tmp674 = (w_sys_tmp675 + r_run_k_20);
	assign w_sys_tmp675 = (r_run_copy3_j_53 * w_sys_tmp668);
	assign w_sys_tmp677 = w_fld_V_3_dataout_1;
	assign w_sys_tmp678 = (w_sys_tmp679 + r_run_k_20);
	assign w_sys_tmp679 = (r_run_copy2_j_52 * w_sys_tmp668);
	assign w_sys_tmp682 = (w_sys_tmp683 + r_run_k_20);
	assign w_sys_tmp683 = (r_run_copy1_j_51 * w_sys_tmp668);
	assign w_sys_tmp685 = w_fld_T_0_dataout_1;
	assign w_sys_tmp686 = (w_sys_tmp687 + r_run_k_20);
	assign w_sys_tmp687 = (r_run_copy0_j_50 * w_sys_tmp668);
	assign w_sys_tmp689 = (r_run_copy0_j_50 + w_sys_intOne);
	assign w_sys_tmp690 = (r_run_copy1_j_51 + w_sys_intOne);
	assign w_sys_tmp691 = (r_run_copy2_j_52 + w_sys_intOne);
	assign w_sys_tmp692 = (r_run_copy3_j_53 + w_sys_intOne);
	assign w_sys_tmp693 = (r_run_copy4_j_54 + w_sys_intOne);
	assign w_sys_tmp694 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp875 = 32'sh00000060;
	assign w_sys_tmp876 = ( !w_sys_tmp877 );
	assign w_sys_tmp877 = (w_sys_tmp878 < r_run_j_21);
	assign w_sys_tmp878 = 32'sh00000081;
	assign w_sys_tmp881 = (w_sys_tmp882 + r_run_k_20);
	assign w_sys_tmp882 = (r_run_j_21 * w_sys_tmp883);
	assign w_sys_tmp883 = 32'sh00000081;
	assign w_sys_tmp884 = w_fld_U_2_dataout_1;
	assign w_sys_tmp885 = (w_sys_tmp886 + r_run_k_20);
	assign w_sys_tmp886 = (r_run_copy4_j_59 * w_sys_tmp883);
	assign w_sys_tmp889 = (w_sys_tmp890 + r_run_k_20);
	assign w_sys_tmp890 = (r_run_copy3_j_58 * w_sys_tmp883);
	assign w_sys_tmp892 = w_fld_V_3_dataout_1;
	assign w_sys_tmp893 = (w_sys_tmp894 + r_run_k_20);
	assign w_sys_tmp894 = (r_run_copy2_j_57 * w_sys_tmp883);
	assign w_sys_tmp897 = (w_sys_tmp898 + r_run_k_20);
	assign w_sys_tmp898 = (r_run_copy1_j_56 * w_sys_tmp883);
	assign w_sys_tmp900 = w_fld_T_0_dataout_1;
	assign w_sys_tmp901 = (w_sys_tmp902 + r_run_k_20);
	assign w_sys_tmp902 = (r_run_copy0_j_55 * w_sys_tmp883);
	assign w_sys_tmp904 = (r_run_copy0_j_55 + w_sys_intOne);
	assign w_sys_tmp905 = (r_run_copy1_j_56 + w_sys_intOne);
	assign w_sys_tmp906 = (r_run_copy2_j_57 + w_sys_intOne);
	assign w_sys_tmp907 = (r_run_copy3_j_58 + w_sys_intOne);
	assign w_sys_tmp908 = (r_run_copy4_j_59 + w_sys_intOne);
	assign w_sys_tmp909 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp1090 = 32'sh00000020;
	assign w_sys_tmp1091 = ( !w_sys_tmp1092 );
	assign w_sys_tmp1092 = (w_sys_tmp1093 < r_run_k_20);
	assign w_sys_tmp1093 = 32'sh00000041;
	assign w_sys_tmp1094 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp1095 = ( !w_sys_tmp1096 );
	assign w_sys_tmp1096 = (w_sys_tmp1097 < r_run_j_21);
	assign w_sys_tmp1097 = 32'sh00000021;
	assign w_sys_tmp1100 = (w_sys_tmp1101 + r_run_k_20);
	assign w_sys_tmp1101 = (r_run_j_21 * w_sys_tmp1102);
	assign w_sys_tmp1102 = 32'sh00000081;
	assign w_sys_tmp1103 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1104 = (w_sys_tmp1105 + r_run_k_20);
	assign w_sys_tmp1105 = (r_run_copy4_j_64 * w_sys_tmp1102);
	assign w_sys_tmp1108 = (w_sys_tmp1109 + r_run_k_20);
	assign w_sys_tmp1109 = (r_run_copy3_j_63 * w_sys_tmp1102);
	assign w_sys_tmp1111 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1112 = (w_sys_tmp1113 + r_run_k_20);
	assign w_sys_tmp1113 = (r_run_copy2_j_62 * w_sys_tmp1102);
	assign w_sys_tmp1116 = (w_sys_tmp1117 + r_run_k_20);
	assign w_sys_tmp1117 = (r_run_copy1_j_61 * w_sys_tmp1102);
	assign w_sys_tmp1119 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1120 = (w_sys_tmp1121 + r_run_k_20);
	assign w_sys_tmp1121 = (r_run_copy0_j_60 * w_sys_tmp1102);
	assign w_sys_tmp1123 = (r_run_copy0_j_60 + w_sys_intOne);
	assign w_sys_tmp1124 = (r_run_copy1_j_61 + w_sys_intOne);
	assign w_sys_tmp1125 = (r_run_copy2_j_62 + w_sys_intOne);
	assign w_sys_tmp1126 = (r_run_copy3_j_63 + w_sys_intOne);
	assign w_sys_tmp1127 = (r_run_copy4_j_64 + w_sys_intOne);
	assign w_sys_tmp1128 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp1309 = 32'sh00000020;
	assign w_sys_tmp1310 = ( !w_sys_tmp1311 );
	assign w_sys_tmp1311 = (w_sys_tmp1312 < r_run_j_21);
	assign w_sys_tmp1312 = 32'sh00000041;
	assign w_sys_tmp1315 = (w_sys_tmp1316 + r_run_k_20);
	assign w_sys_tmp1316 = (r_run_j_21 * w_sys_tmp1317);
	assign w_sys_tmp1317 = 32'sh00000081;
	assign w_sys_tmp1318 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1319 = (w_sys_tmp1320 + r_run_k_20);
	assign w_sys_tmp1320 = (r_run_copy4_j_69 * w_sys_tmp1317);
	assign w_sys_tmp1323 = (w_sys_tmp1324 + r_run_k_20);
	assign w_sys_tmp1324 = (r_run_copy3_j_68 * w_sys_tmp1317);
	assign w_sys_tmp1326 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1327 = (w_sys_tmp1328 + r_run_k_20);
	assign w_sys_tmp1328 = (r_run_copy2_j_67 * w_sys_tmp1317);
	assign w_sys_tmp1331 = (w_sys_tmp1332 + r_run_k_20);
	assign w_sys_tmp1332 = (r_run_copy1_j_66 * w_sys_tmp1317);
	assign w_sys_tmp1334 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1335 = (w_sys_tmp1336 + r_run_k_20);
	assign w_sys_tmp1336 = (r_run_copy0_j_65 * w_sys_tmp1317);
	assign w_sys_tmp1338 = (r_run_copy0_j_65 + w_sys_intOne);
	assign w_sys_tmp1339 = (r_run_copy1_j_66 + w_sys_intOne);
	assign w_sys_tmp1340 = (r_run_copy2_j_67 + w_sys_intOne);
	assign w_sys_tmp1341 = (r_run_copy3_j_68 + w_sys_intOne);
	assign w_sys_tmp1342 = (r_run_copy4_j_69 + w_sys_intOne);
	assign w_sys_tmp1343 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp1524 = 32'sh00000040;
	assign w_sys_tmp1525 = ( !w_sys_tmp1526 );
	assign w_sys_tmp1526 = (w_sys_tmp1527 < r_run_j_21);
	assign w_sys_tmp1527 = 32'sh00000061;
	assign w_sys_tmp1530 = (w_sys_tmp1531 + r_run_k_20);
	assign w_sys_tmp1531 = (r_run_j_21 * w_sys_tmp1532);
	assign w_sys_tmp1532 = 32'sh00000081;
	assign w_sys_tmp1533 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1534 = (w_sys_tmp1535 + r_run_k_20);
	assign w_sys_tmp1535 = (r_run_copy4_j_74 * w_sys_tmp1532);
	assign w_sys_tmp1538 = (w_sys_tmp1539 + r_run_k_20);
	assign w_sys_tmp1539 = (r_run_copy3_j_73 * w_sys_tmp1532);
	assign w_sys_tmp1541 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1542 = (w_sys_tmp1543 + r_run_k_20);
	assign w_sys_tmp1543 = (r_run_copy2_j_72 * w_sys_tmp1532);
	assign w_sys_tmp1546 = (w_sys_tmp1547 + r_run_k_20);
	assign w_sys_tmp1547 = (r_run_copy1_j_71 * w_sys_tmp1532);
	assign w_sys_tmp1549 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1550 = (w_sys_tmp1551 + r_run_k_20);
	assign w_sys_tmp1551 = (r_run_copy0_j_70 * w_sys_tmp1532);
	assign w_sys_tmp1553 = (r_run_copy0_j_70 + w_sys_intOne);
	assign w_sys_tmp1554 = (r_run_copy1_j_71 + w_sys_intOne);
	assign w_sys_tmp1555 = (r_run_copy2_j_72 + w_sys_intOne);
	assign w_sys_tmp1556 = (r_run_copy3_j_73 + w_sys_intOne);
	assign w_sys_tmp1557 = (r_run_copy4_j_74 + w_sys_intOne);
	assign w_sys_tmp1558 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp1739 = 32'sh00000060;
	assign w_sys_tmp1740 = ( !w_sys_tmp1741 );
	assign w_sys_tmp1741 = (w_sys_tmp1742 < r_run_j_21);
	assign w_sys_tmp1742 = 32'sh00000081;
	assign w_sys_tmp1745 = (w_sys_tmp1746 + r_run_k_20);
	assign w_sys_tmp1746 = (r_run_j_21 * w_sys_tmp1747);
	assign w_sys_tmp1747 = 32'sh00000081;
	assign w_sys_tmp1748 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1749 = (w_sys_tmp1750 + r_run_k_20);
	assign w_sys_tmp1750 = (r_run_copy4_j_79 * w_sys_tmp1747);
	assign w_sys_tmp1753 = (w_sys_tmp1754 + r_run_k_20);
	assign w_sys_tmp1754 = (r_run_copy3_j_78 * w_sys_tmp1747);
	assign w_sys_tmp1756 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1757 = (w_sys_tmp1758 + r_run_k_20);
	assign w_sys_tmp1758 = (r_run_copy2_j_77 * w_sys_tmp1747);
	assign w_sys_tmp1761 = (w_sys_tmp1762 + r_run_k_20);
	assign w_sys_tmp1762 = (r_run_copy1_j_76 * w_sys_tmp1747);
	assign w_sys_tmp1764 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1765 = (w_sys_tmp1766 + r_run_k_20);
	assign w_sys_tmp1766 = (r_run_copy0_j_75 * w_sys_tmp1747);
	assign w_sys_tmp1768 = (r_run_copy0_j_75 + w_sys_intOne);
	assign w_sys_tmp1769 = (r_run_copy1_j_76 + w_sys_intOne);
	assign w_sys_tmp1770 = (r_run_copy2_j_77 + w_sys_intOne);
	assign w_sys_tmp1771 = (r_run_copy3_j_78 + w_sys_intOne);
	assign w_sys_tmp1772 = (r_run_copy4_j_79 + w_sys_intOne);
	assign w_sys_tmp1773 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp1954 = 32'sh00000040;
	assign w_sys_tmp1955 = ( !w_sys_tmp1956 );
	assign w_sys_tmp1956 = (w_sys_tmp1957 < r_run_k_20);
	assign w_sys_tmp1957 = 32'sh00000061;
	assign w_sys_tmp1958 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp1959 = ( !w_sys_tmp1960 );
	assign w_sys_tmp1960 = (w_sys_tmp1961 < r_run_j_21);
	assign w_sys_tmp1961 = 32'sh00000021;
	assign w_sys_tmp1964 = (w_sys_tmp1965 + r_run_k_20);
	assign w_sys_tmp1965 = (r_run_j_21 * w_sys_tmp1966);
	assign w_sys_tmp1966 = 32'sh00000081;
	assign w_sys_tmp1967 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1968 = (w_sys_tmp1969 + r_run_k_20);
	assign w_sys_tmp1969 = (r_run_copy4_j_84 * w_sys_tmp1966);
	assign w_sys_tmp1972 = (w_sys_tmp1973 + r_run_k_20);
	assign w_sys_tmp1973 = (r_run_copy3_j_83 * w_sys_tmp1966);
	assign w_sys_tmp1975 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1976 = (w_sys_tmp1977 + r_run_k_20);
	assign w_sys_tmp1977 = (r_run_copy2_j_82 * w_sys_tmp1966);
	assign w_sys_tmp1980 = (w_sys_tmp1981 + r_run_k_20);
	assign w_sys_tmp1981 = (r_run_copy1_j_81 * w_sys_tmp1966);
	assign w_sys_tmp1983 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1984 = (w_sys_tmp1985 + r_run_k_20);
	assign w_sys_tmp1985 = (r_run_copy0_j_80 * w_sys_tmp1966);
	assign w_sys_tmp1987 = (r_run_copy0_j_80 + w_sys_intOne);
	assign w_sys_tmp1988 = (r_run_copy1_j_81 + w_sys_intOne);
	assign w_sys_tmp1989 = (r_run_copy2_j_82 + w_sys_intOne);
	assign w_sys_tmp1990 = (r_run_copy3_j_83 + w_sys_intOne);
	assign w_sys_tmp1991 = (r_run_copy4_j_84 + w_sys_intOne);
	assign w_sys_tmp1992 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp2173 = 32'sh00000020;
	assign w_sys_tmp2174 = ( !w_sys_tmp2175 );
	assign w_sys_tmp2175 = (w_sys_tmp2176 < r_run_j_21);
	assign w_sys_tmp2176 = 32'sh00000041;
	assign w_sys_tmp2179 = (w_sys_tmp2180 + r_run_k_20);
	assign w_sys_tmp2180 = (r_run_j_21 * w_sys_tmp2181);
	assign w_sys_tmp2181 = 32'sh00000081;
	assign w_sys_tmp2182 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2183 = (w_sys_tmp2184 + r_run_k_20);
	assign w_sys_tmp2184 = (r_run_copy4_j_89 * w_sys_tmp2181);
	assign w_sys_tmp2187 = (w_sys_tmp2188 + r_run_k_20);
	assign w_sys_tmp2188 = (r_run_copy3_j_88 * w_sys_tmp2181);
	assign w_sys_tmp2190 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2191 = (w_sys_tmp2192 + r_run_k_20);
	assign w_sys_tmp2192 = (r_run_copy2_j_87 * w_sys_tmp2181);
	assign w_sys_tmp2195 = (w_sys_tmp2196 + r_run_k_20);
	assign w_sys_tmp2196 = (r_run_copy1_j_86 * w_sys_tmp2181);
	assign w_sys_tmp2198 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2199 = (w_sys_tmp2200 + r_run_k_20);
	assign w_sys_tmp2200 = (r_run_copy0_j_85 * w_sys_tmp2181);
	assign w_sys_tmp2202 = (r_run_copy0_j_85 + w_sys_intOne);
	assign w_sys_tmp2203 = (r_run_copy1_j_86 + w_sys_intOne);
	assign w_sys_tmp2204 = (r_run_copy2_j_87 + w_sys_intOne);
	assign w_sys_tmp2205 = (r_run_copy3_j_88 + w_sys_intOne);
	assign w_sys_tmp2206 = (r_run_copy4_j_89 + w_sys_intOne);
	assign w_sys_tmp2207 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp2388 = 32'sh00000040;
	assign w_sys_tmp2389 = ( !w_sys_tmp2390 );
	assign w_sys_tmp2390 = (w_sys_tmp2391 < r_run_j_21);
	assign w_sys_tmp2391 = 32'sh00000061;
	assign w_sys_tmp2394 = (w_sys_tmp2395 + r_run_k_20);
	assign w_sys_tmp2395 = (r_run_j_21 * w_sys_tmp2396);
	assign w_sys_tmp2396 = 32'sh00000081;
	assign w_sys_tmp2397 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2398 = (w_sys_tmp2399 + r_run_k_20);
	assign w_sys_tmp2399 = (r_run_copy4_j_94 * w_sys_tmp2396);
	assign w_sys_tmp2402 = (w_sys_tmp2403 + r_run_k_20);
	assign w_sys_tmp2403 = (r_run_copy3_j_93 * w_sys_tmp2396);
	assign w_sys_tmp2405 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2406 = (w_sys_tmp2407 + r_run_k_20);
	assign w_sys_tmp2407 = (r_run_copy2_j_92 * w_sys_tmp2396);
	assign w_sys_tmp2410 = (w_sys_tmp2411 + r_run_k_20);
	assign w_sys_tmp2411 = (r_run_copy1_j_91 * w_sys_tmp2396);
	assign w_sys_tmp2413 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2414 = (w_sys_tmp2415 + r_run_k_20);
	assign w_sys_tmp2415 = (r_run_copy0_j_90 * w_sys_tmp2396);
	assign w_sys_tmp2417 = (r_run_copy0_j_90 + w_sys_intOne);
	assign w_sys_tmp2418 = (r_run_copy1_j_91 + w_sys_intOne);
	assign w_sys_tmp2419 = (r_run_copy2_j_92 + w_sys_intOne);
	assign w_sys_tmp2420 = (r_run_copy3_j_93 + w_sys_intOne);
	assign w_sys_tmp2421 = (r_run_copy4_j_94 + w_sys_intOne);
	assign w_sys_tmp2422 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp2603 = 32'sh00000060;
	assign w_sys_tmp2604 = ( !w_sys_tmp2605 );
	assign w_sys_tmp2605 = (w_sys_tmp2606 < r_run_j_21);
	assign w_sys_tmp2606 = 32'sh00000081;
	assign w_sys_tmp2609 = (w_sys_tmp2610 + r_run_k_20);
	assign w_sys_tmp2610 = (r_run_j_21 * w_sys_tmp2611);
	assign w_sys_tmp2611 = 32'sh00000081;
	assign w_sys_tmp2612 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2613 = (w_sys_tmp2614 + r_run_k_20);
	assign w_sys_tmp2614 = (r_run_copy4_j_99 * w_sys_tmp2611);
	assign w_sys_tmp2617 = (w_sys_tmp2618 + r_run_k_20);
	assign w_sys_tmp2618 = (r_run_copy3_j_98 * w_sys_tmp2611);
	assign w_sys_tmp2620 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2621 = (w_sys_tmp2622 + r_run_k_20);
	assign w_sys_tmp2622 = (r_run_copy2_j_97 * w_sys_tmp2611);
	assign w_sys_tmp2625 = (w_sys_tmp2626 + r_run_k_20);
	assign w_sys_tmp2626 = (r_run_copy1_j_96 * w_sys_tmp2611);
	assign w_sys_tmp2628 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2629 = (w_sys_tmp2630 + r_run_k_20);
	assign w_sys_tmp2630 = (r_run_copy0_j_95 * w_sys_tmp2611);
	assign w_sys_tmp2632 = (r_run_copy0_j_95 + w_sys_intOne);
	assign w_sys_tmp2633 = (r_run_copy1_j_96 + w_sys_intOne);
	assign w_sys_tmp2634 = (r_run_copy2_j_97 + w_sys_intOne);
	assign w_sys_tmp2635 = (r_run_copy3_j_98 + w_sys_intOne);
	assign w_sys_tmp2636 = (r_run_copy4_j_99 + w_sys_intOne);
	assign w_sys_tmp2637 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp2818 = 32'sh00000060;
	assign w_sys_tmp2819 = ( !w_sys_tmp2820 );
	assign w_sys_tmp2820 = (w_sys_tmp2821 < r_run_k_20);
	assign w_sys_tmp2821 = 32'sh00000081;
	assign w_sys_tmp2822 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp2823 = ( !w_sys_tmp2824 );
	assign w_sys_tmp2824 = (w_sys_tmp2825 < r_run_j_21);
	assign w_sys_tmp2825 = 32'sh00000021;
	assign w_sys_tmp2828 = (w_sys_tmp2829 + r_run_k_20);
	assign w_sys_tmp2829 = (r_run_j_21 * w_sys_tmp2830);
	assign w_sys_tmp2830 = 32'sh00000081;
	assign w_sys_tmp2831 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2832 = (w_sys_tmp2833 + r_run_k_20);
	assign w_sys_tmp2833 = (r_run_copy4_j_104 * w_sys_tmp2830);
	assign w_sys_tmp2836 = (w_sys_tmp2837 + r_run_k_20);
	assign w_sys_tmp2837 = (r_run_copy3_j_103 * w_sys_tmp2830);
	assign w_sys_tmp2839 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2840 = (w_sys_tmp2841 + r_run_k_20);
	assign w_sys_tmp2841 = (r_run_copy2_j_102 * w_sys_tmp2830);
	assign w_sys_tmp2844 = (w_sys_tmp2845 + r_run_k_20);
	assign w_sys_tmp2845 = (r_run_copy1_j_101 * w_sys_tmp2830);
	assign w_sys_tmp2847 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2848 = (w_sys_tmp2849 + r_run_k_20);
	assign w_sys_tmp2849 = (r_run_copy0_j_100 * w_sys_tmp2830);
	assign w_sys_tmp2851 = (r_run_copy0_j_100 + w_sys_intOne);
	assign w_sys_tmp2852 = (r_run_copy1_j_101 + w_sys_intOne);
	assign w_sys_tmp2853 = (r_run_copy2_j_102 + w_sys_intOne);
	assign w_sys_tmp2854 = (r_run_copy3_j_103 + w_sys_intOne);
	assign w_sys_tmp2855 = (r_run_copy4_j_104 + w_sys_intOne);
	assign w_sys_tmp2856 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp3037 = 32'sh00000020;
	assign w_sys_tmp3038 = ( !w_sys_tmp3039 );
	assign w_sys_tmp3039 = (w_sys_tmp3040 < r_run_j_21);
	assign w_sys_tmp3040 = 32'sh00000041;
	assign w_sys_tmp3043 = (w_sys_tmp3044 + r_run_k_20);
	assign w_sys_tmp3044 = (r_run_j_21 * w_sys_tmp3045);
	assign w_sys_tmp3045 = 32'sh00000081;
	assign w_sys_tmp3046 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3047 = (w_sys_tmp3048 + r_run_k_20);
	assign w_sys_tmp3048 = (r_run_copy4_j_109 * w_sys_tmp3045);
	assign w_sys_tmp3051 = (w_sys_tmp3052 + r_run_k_20);
	assign w_sys_tmp3052 = (r_run_copy3_j_108 * w_sys_tmp3045);
	assign w_sys_tmp3054 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3055 = (w_sys_tmp3056 + r_run_k_20);
	assign w_sys_tmp3056 = (r_run_copy2_j_107 * w_sys_tmp3045);
	assign w_sys_tmp3059 = (w_sys_tmp3060 + r_run_k_20);
	assign w_sys_tmp3060 = (r_run_copy1_j_106 * w_sys_tmp3045);
	assign w_sys_tmp3062 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3063 = (w_sys_tmp3064 + r_run_k_20);
	assign w_sys_tmp3064 = (r_run_copy0_j_105 * w_sys_tmp3045);
	assign w_sys_tmp3066 = (r_run_copy0_j_105 + w_sys_intOne);
	assign w_sys_tmp3067 = (r_run_copy1_j_106 + w_sys_intOne);
	assign w_sys_tmp3068 = (r_run_copy2_j_107 + w_sys_intOne);
	assign w_sys_tmp3069 = (r_run_copy3_j_108 + w_sys_intOne);
	assign w_sys_tmp3070 = (r_run_copy4_j_109 + w_sys_intOne);
	assign w_sys_tmp3071 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp3252 = 32'sh00000040;
	assign w_sys_tmp3253 = ( !w_sys_tmp3254 );
	assign w_sys_tmp3254 = (w_sys_tmp3255 < r_run_j_21);
	assign w_sys_tmp3255 = 32'sh00000061;
	assign w_sys_tmp3258 = (w_sys_tmp3259 + r_run_k_20);
	assign w_sys_tmp3259 = (r_run_j_21 * w_sys_tmp3260);
	assign w_sys_tmp3260 = 32'sh00000081;
	assign w_sys_tmp3261 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3262 = (w_sys_tmp3263 + r_run_k_20);
	assign w_sys_tmp3263 = (r_run_copy4_j_114 * w_sys_tmp3260);
	assign w_sys_tmp3266 = (w_sys_tmp3267 + r_run_k_20);
	assign w_sys_tmp3267 = (r_run_copy3_j_113 * w_sys_tmp3260);
	assign w_sys_tmp3269 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3270 = (w_sys_tmp3271 + r_run_k_20);
	assign w_sys_tmp3271 = (r_run_copy2_j_112 * w_sys_tmp3260);
	assign w_sys_tmp3274 = (w_sys_tmp3275 + r_run_k_20);
	assign w_sys_tmp3275 = (r_run_copy1_j_111 * w_sys_tmp3260);
	assign w_sys_tmp3277 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3278 = (w_sys_tmp3279 + r_run_k_20);
	assign w_sys_tmp3279 = (r_run_copy0_j_110 * w_sys_tmp3260);
	assign w_sys_tmp3281 = (r_run_copy0_j_110 + w_sys_intOne);
	assign w_sys_tmp3282 = (r_run_copy1_j_111 + w_sys_intOne);
	assign w_sys_tmp3283 = (r_run_copy2_j_112 + w_sys_intOne);
	assign w_sys_tmp3284 = (r_run_copy3_j_113 + w_sys_intOne);
	assign w_sys_tmp3285 = (r_run_copy4_j_114 + w_sys_intOne);
	assign w_sys_tmp3286 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp3467 = 32'sh00000060;
	assign w_sys_tmp3468 = ( !w_sys_tmp3469 );
	assign w_sys_tmp3469 = (w_sys_tmp3470 < r_run_j_21);
	assign w_sys_tmp3470 = 32'sh00000081;
	assign w_sys_tmp3473 = (w_sys_tmp3474 + r_run_k_20);
	assign w_sys_tmp3474 = (r_run_j_21 * w_sys_tmp3475);
	assign w_sys_tmp3475 = 32'sh00000081;
	assign w_sys_tmp3476 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3477 = (w_sys_tmp3478 + r_run_k_20);
	assign w_sys_tmp3478 = (r_run_copy4_j_119 * w_sys_tmp3475);
	assign w_sys_tmp3481 = (w_sys_tmp3482 + r_run_k_20);
	assign w_sys_tmp3482 = (r_run_copy3_j_118 * w_sys_tmp3475);
	assign w_sys_tmp3484 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3485 = (w_sys_tmp3486 + r_run_k_20);
	assign w_sys_tmp3486 = (r_run_copy2_j_117 * w_sys_tmp3475);
	assign w_sys_tmp3489 = (w_sys_tmp3490 + r_run_k_20);
	assign w_sys_tmp3490 = (r_run_copy1_j_116 * w_sys_tmp3475);
	assign w_sys_tmp3492 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3493 = (w_sys_tmp3494 + r_run_k_20);
	assign w_sys_tmp3494 = (r_run_copy0_j_115 * w_sys_tmp3475);
	assign w_sys_tmp3496 = (r_run_copy0_j_115 + w_sys_intOne);
	assign w_sys_tmp3497 = (r_run_copy1_j_116 + w_sys_intOne);
	assign w_sys_tmp3498 = (r_run_copy2_j_117 + w_sys_intOne);
	assign w_sys_tmp3499 = (r_run_copy3_j_118 + w_sys_intOne);
	assign w_sys_tmp3500 = (r_run_copy4_j_119 + w_sys_intOne);
	assign w_sys_tmp3501 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp3682 = ( !w_sys_tmp3683 );
	assign w_sys_tmp3683 = (r_run_nlast_35 < r_run_n_22);
	assign w_sys_tmp3684 = (r_run_n_22 + w_sys_intOne);
	assign w_sys_tmp3685 = 32'sh00000002;
	assign w_sys_tmp3686 = ( !w_sys_tmp3687 );
	assign w_sys_tmp3687 = (w_sys_tmp3688 < r_run_k_20);
	assign w_sys_tmp3688 = 32'sh00000020;
	assign w_sys_tmp3691 = (w_sys_tmp3692 + r_run_k_20);
	assign w_sys_tmp3692 = 32'sh000010a1;
	assign w_sys_tmp3693 = w_sub01_result_dataout;
	assign w_sys_tmp3694 = (w_sys_tmp3695 + r_run_k_20);
	assign w_sys_tmp3695 = 32'sh00000102;
	assign w_sys_tmp3697 = (w_sys_tmp3698 + r_run_k_20);
	assign w_sys_tmp3698 = 32'sh00000081;
	assign w_sys_tmp3699 = w_sub00_result_dataout;
	assign w_sys_tmp3700 = (w_sys_tmp3701 + r_run_k_20);
	assign w_sys_tmp3701 = 32'sh00001020;
	assign w_sys_tmp3703 = (w_sys_tmp3704 + r_run_k_20);
	assign w_sys_tmp3704 = 32'sh00001122;
	assign w_sys_tmp3721 = w_sub02_result_dataout;
	assign w_sys_tmp3724 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp3725 = 32'sh00000021;
	assign w_sys_tmp3726 = ( !w_sys_tmp3727 );
	assign w_sys_tmp3727 = (w_sys_tmp3728 < r_run_k_20);
	assign w_sys_tmp3728 = 32'sh00000040;
	assign w_sys_tmp3731 = (w_sys_tmp3732 + r_run_k_20);
	assign w_sys_tmp3732 = 32'sh000010a1;
	assign w_sys_tmp3733 = w_sub05_result_dataout;
	assign w_sys_tmp3734 = (w_sys_tmp3735 + r_run_k_20);
	assign w_sys_tmp3735 = 32'sh00000102;
	assign w_sys_tmp3737 = (w_sys_tmp3738 + r_run_k_20);
	assign w_sys_tmp3738 = 32'sh00000081;
	assign w_sys_tmp3739 = w_sub04_result_dataout;
	assign w_sys_tmp3740 = (w_sys_tmp3741 + r_run_k_20);
	assign w_sys_tmp3741 = 32'sh00001020;
	assign w_sys_tmp3743 = (w_sys_tmp3744 + r_run_k_20);
	assign w_sys_tmp3744 = 32'sh00001122;
	assign w_sys_tmp3761 = w_sub06_result_dataout;
	assign w_sys_tmp3764 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp3765 = 32'sh00000041;
	assign w_sys_tmp3766 = ( !w_sys_tmp3767 );
	assign w_sys_tmp3767 = (w_sys_tmp3768 < r_run_k_20);
	assign w_sys_tmp3768 = 32'sh00000060;
	assign w_sys_tmp3771 = (w_sys_tmp3772 + r_run_k_20);
	assign w_sys_tmp3772 = 32'sh000010a1;
	assign w_sys_tmp3773 = w_sub09_result_dataout;
	assign w_sys_tmp3774 = (w_sys_tmp3775 + r_run_k_20);
	assign w_sys_tmp3775 = 32'sh00000102;
	assign w_sys_tmp3777 = (w_sys_tmp3778 + r_run_k_20);
	assign w_sys_tmp3778 = 32'sh00000081;
	assign w_sys_tmp3779 = w_sub08_result_dataout;
	assign w_sys_tmp3780 = (w_sys_tmp3781 + r_run_k_20);
	assign w_sys_tmp3781 = 32'sh00001020;
	assign w_sys_tmp3783 = (w_sys_tmp3784 + r_run_k_20);
	assign w_sys_tmp3784 = 32'sh00001122;
	assign w_sys_tmp3801 = w_sub10_result_dataout;
	assign w_sys_tmp3804 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp3805 = 32'sh00000061;
	assign w_sys_tmp3806 = ( !w_sys_tmp3807 );
	assign w_sys_tmp3807 = (w_sys_tmp3808 < r_run_k_20);
	assign w_sys_tmp3808 = 32'sh00000080;
	assign w_sys_tmp3811 = (w_sys_tmp3812 + r_run_k_20);
	assign w_sys_tmp3812 = 32'sh000010a1;
	assign w_sys_tmp3813 = w_sub13_result_dataout;
	assign w_sys_tmp3814 = (w_sys_tmp3815 + r_run_k_20);
	assign w_sys_tmp3815 = 32'sh00000102;
	assign w_sys_tmp3817 = (w_sys_tmp3818 + r_run_k_20);
	assign w_sys_tmp3818 = 32'sh00000081;
	assign w_sys_tmp3819 = w_sub12_result_dataout;
	assign w_sys_tmp3820 = (w_sys_tmp3821 + r_run_k_20);
	assign w_sys_tmp3821 = 32'sh00001020;
	assign w_sys_tmp3823 = (w_sys_tmp3824 + r_run_k_20);
	assign w_sys_tmp3824 = 32'sh00001122;
	assign w_sys_tmp3841 = w_sub14_result_dataout;
	assign w_sys_tmp3842 = (w_sys_tmp3843 + r_run_k_20);
	assign w_sys_tmp3843 = 32'sh00000183;
	assign w_sys_tmp3844 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp3845 = 32'sh00000002;
	assign w_sys_tmp3846 = ( !w_sys_tmp3847 );
	assign w_sys_tmp3847 = (w_sys_tmp3848 < r_run_j_21);
	assign w_sys_tmp3848 = 32'sh00000020;
	assign w_sys_tmp3851 = (w_sys_tmp3852 + w_sys_tmp3854);
	assign w_sys_tmp3852 = (r_run_j_21 * w_sys_tmp3853);
	assign w_sys_tmp3853 = 32'sh00000081;
	assign w_sys_tmp3854 = 32'sh00000021;
	assign w_sys_tmp3855 = w_sub04_result_dataout;
	assign w_sys_tmp3856 = (w_sys_tmp3857 + w_sys_tmp3854);
	assign w_sys_tmp3857 = (r_run_copy10_j_130 * w_sys_tmp3853);
	assign w_sys_tmp3861 = (w_sys_tmp3862 + w_sys_tmp3864);
	assign w_sys_tmp3862 = (r_run_copy9_j_129 * w_sys_tmp3853);
	assign w_sys_tmp3864 = 32'sh00000020;
	assign w_sys_tmp3865 = w_sub00_result_dataout;
	assign w_sys_tmp3866 = (w_sys_tmp3867 + w_sys_tmp3864);
	assign w_sys_tmp3867 = (r_run_copy8_j_128 * w_sys_tmp3853);
	assign w_sys_tmp3871 = (w_sys_tmp3872 + w_sys_tmp3874);
	assign w_sys_tmp3872 = (r_run_copy7_j_127 * w_sys_tmp3853);
	assign w_sys_tmp3874 = 32'sh00000041;
	assign w_sys_tmp3875 = (w_sys_tmp3876 + w_sys_tmp3874);
	assign w_sys_tmp3876 = (r_run_copy6_j_126 * w_sys_tmp3853);
	assign w_sys_tmp3880 = (w_sys_tmp3881 + w_sys_tmp3883);
	assign w_sys_tmp3881 = (r_run_copy5_j_125 * w_sys_tmp3853);
	assign w_sys_tmp3883 = 32'sh00000040;
	assign w_sys_tmp3885 = (w_sys_tmp3886 + w_sys_tmp3883);
	assign w_sys_tmp3886 = (r_run_copy4_j_124 * w_sys_tmp3853);
	assign w_sys_tmp3890 = (w_sys_tmp3891 + w_sys_tmp3893);
	assign w_sys_tmp3891 = (r_run_copy3_j_123 * w_sys_tmp3853);
	assign w_sys_tmp3893 = 32'sh00000061;
	assign w_sys_tmp3894 = (w_sys_tmp3895 + w_sys_tmp3893);
	assign w_sys_tmp3895 = (r_run_copy2_j_122 * w_sys_tmp3853);
	assign w_sys_tmp3899 = (w_sys_tmp3900 + w_sys_tmp3902);
	assign w_sys_tmp3900 = (r_run_copy1_j_121 * w_sys_tmp3853);
	assign w_sys_tmp3902 = 32'sh00000060;
	assign w_sys_tmp3903 = w_sub08_result_dataout;
	assign w_sys_tmp3904 = (w_sys_tmp3905 + w_sys_tmp3902);
	assign w_sys_tmp3905 = (r_run_copy0_j_120 * w_sys_tmp3853);
	assign w_sys_tmp3908 = (r_run_copy0_j_120 + w_sys_intOne);
	assign w_sys_tmp3909 = (r_run_copy1_j_121 + w_sys_intOne);
	assign w_sys_tmp3910 = (r_run_copy2_j_122 + w_sys_intOne);
	assign w_sys_tmp3911 = (r_run_copy3_j_123 + w_sys_intOne);
	assign w_sys_tmp3912 = (r_run_copy4_j_124 + w_sys_intOne);
	assign w_sys_tmp3913 = (r_run_copy5_j_125 + w_sys_intOne);
	assign w_sys_tmp3914 = (r_run_copy6_j_126 + w_sys_intOne);
	assign w_sys_tmp3915 = (r_run_copy7_j_127 + w_sys_intOne);
	assign w_sys_tmp3916 = (r_run_copy8_j_128 + w_sys_intOne);
	assign w_sys_tmp3917 = (r_run_copy9_j_129 + w_sys_intOne);
	assign w_sys_tmp3918 = (r_run_copy10_j_130 + w_sys_intOne);
	assign w_sys_tmp3919 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp4346 = 32'sh00000021;
	assign w_sys_tmp4347 = ( !w_sys_tmp4348 );
	assign w_sys_tmp4348 = (w_sys_tmp4349 < r_run_j_21);
	assign w_sys_tmp4349 = 32'sh00000040;
	assign w_sys_tmp4351 = (r_run_j_21 - w_sys_tmp4352);
	assign w_sys_tmp4352 = 32'sh0000001f;
	assign w_sys_tmp4354 = (w_sys_tmp4355 + w_sys_tmp4357);
	assign w_sys_tmp4355 = (r_run_tmpj_36 * w_sys_tmp4356);
	assign w_sys_tmp4356 = 32'sh00000081;
	assign w_sys_tmp4357 = 32'sh00000021;
	assign w_sys_tmp4358 = w_sub05_result_dataout;
	assign w_sys_tmp4359 = (w_sys_tmp4360 + w_sys_tmp4357);
	assign w_sys_tmp4360 = (w_sys_tmp4361 * w_sys_tmp4356);
	assign w_sys_tmp4361 = w_sys_tmp4351;
	assign w_sys_tmp4365 = (w_sys_tmp4355 + w_sys_tmp4368);
	assign w_sys_tmp4368 = 32'sh00000020;
	assign w_sys_tmp4369 = w_sub01_result_dataout;
	assign w_sys_tmp4375 = (w_sys_tmp4355 + w_sys_tmp4378);
	assign w_sys_tmp4378 = 32'sh00000041;
	assign w_sys_tmp4379 = (w_sys_tmp4360 + w_sys_tmp4378);
	assign w_sys_tmp4385 = (w_sys_tmp4355 + w_sys_tmp4388);
	assign w_sys_tmp4388 = 32'sh00000040;
	assign w_sys_tmp4395 = (w_sys_tmp4355 + w_sys_tmp4398);
	assign w_sys_tmp4398 = 32'sh00000061;
	assign w_sys_tmp4399 = (w_sys_tmp4360 + w_sys_tmp4398);
	assign w_sys_tmp4405 = (w_sys_tmp4355 + w_sys_tmp4408);
	assign w_sys_tmp4408 = 32'sh00000060;
	assign w_sys_tmp4409 = w_sub09_result_dataout;
	assign w_sys_tmp4414 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp4793 = 32'sh00000041;
	assign w_sys_tmp4794 = ( !w_sys_tmp4795 );
	assign w_sys_tmp4795 = (w_sys_tmp4796 < r_run_j_21);
	assign w_sys_tmp4796 = 32'sh00000060;
	assign w_sys_tmp4798 = (r_run_j_21 - w_sys_tmp4799);
	assign w_sys_tmp4799 = 32'sh0000003f;
	assign w_sys_tmp4801 = (w_sys_tmp4802 + w_sys_tmp4804);
	assign w_sys_tmp4802 = (r_run_tmpj_36 * w_sys_tmp4803);
	assign w_sys_tmp4803 = 32'sh00000081;
	assign w_sys_tmp4804 = 32'sh00000021;
	assign w_sys_tmp4805 = w_sub06_result_dataout;
	assign w_sys_tmp4806 = (w_sys_tmp4807 + w_sys_tmp4804);
	assign w_sys_tmp4807 = (w_sys_tmp4808 * w_sys_tmp4803);
	assign w_sys_tmp4808 = w_sys_tmp4798;
	assign w_sys_tmp4812 = (w_sys_tmp4802 + w_sys_tmp4815);
	assign w_sys_tmp4815 = 32'sh00000020;
	assign w_sys_tmp4816 = w_sub02_result_dataout;
	assign w_sys_tmp4822 = (w_sys_tmp4802 + w_sys_tmp4825);
	assign w_sys_tmp4825 = 32'sh00000041;
	assign w_sys_tmp4826 = (w_sys_tmp4807 + w_sys_tmp4825);
	assign w_sys_tmp4832 = (w_sys_tmp4802 + w_sys_tmp4835);
	assign w_sys_tmp4835 = 32'sh00000040;
	assign w_sys_tmp4842 = (w_sys_tmp4802 + w_sys_tmp4845);
	assign w_sys_tmp4845 = 32'sh00000061;
	assign w_sys_tmp4846 = (w_sys_tmp4807 + w_sys_tmp4845);
	assign w_sys_tmp4852 = (w_sys_tmp4802 + w_sys_tmp4855);
	assign w_sys_tmp4855 = 32'sh00000060;
	assign w_sys_tmp4856 = w_sub10_result_dataout;
	assign w_sys_tmp4861 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp5240 = 32'sh00000061;
	assign w_sys_tmp5241 = ( !w_sys_tmp5242 );
	assign w_sys_tmp5242 = (w_sys_tmp5243 < r_run_j_21);
	assign w_sys_tmp5243 = 32'sh00000080;
	assign w_sys_tmp5245 = (r_run_j_21 - w_sys_tmp5246);
	assign w_sys_tmp5246 = 32'sh0000005f;
	assign w_sys_tmp5248 = (w_sys_tmp5249 + w_sys_tmp5251);
	assign w_sys_tmp5249 = (r_run_tmpj_36 * w_sys_tmp5250);
	assign w_sys_tmp5250 = 32'sh00000081;
	assign w_sys_tmp5251 = 32'sh00000021;
	assign w_sys_tmp5252 = w_sub07_result_dataout;
	assign w_sys_tmp5253 = (w_sys_tmp5254 + w_sys_tmp5251);
	assign w_sys_tmp5254 = (w_sys_tmp5255 * w_sys_tmp5250);
	assign w_sys_tmp5255 = w_sys_tmp5245;
	assign w_sys_tmp5259 = (w_sys_tmp5249 + w_sys_tmp5262);
	assign w_sys_tmp5262 = 32'sh00000020;
	assign w_sys_tmp5263 = w_sub03_result_dataout;
	assign w_sys_tmp5269 = (w_sys_tmp5249 + w_sys_tmp5272);
	assign w_sys_tmp5272 = 32'sh00000041;
	assign w_sys_tmp5273 = (w_sys_tmp5254 + w_sys_tmp5272);
	assign w_sys_tmp5279 = (w_sys_tmp5249 + w_sys_tmp5282);
	assign w_sys_tmp5282 = 32'sh00000040;
	assign w_sys_tmp5289 = (w_sys_tmp5249 + w_sys_tmp5292);
	assign w_sys_tmp5292 = 32'sh00000061;
	assign w_sys_tmp5293 = (w_sys_tmp5254 + w_sys_tmp5292);
	assign w_sys_tmp5299 = (w_sys_tmp5249 + w_sys_tmp5302);
	assign w_sys_tmp5302 = 32'sh00000060;
	assign w_sys_tmp5303 = w_sub11_result_dataout;
	assign w_sys_tmp5308 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp5687 = 32'sh00000002;
	assign w_sys_tmp5688 = ( !w_sys_tmp5689 );
	assign w_sys_tmp5689 = (w_sys_tmp5690 < r_run_k_20);
	assign w_sys_tmp5690 = 32'sh00000020;
	assign w_sys_tmp5691 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp5692 = 32'sh00000002;
	assign w_sys_tmp5693 = ( !w_sys_tmp5694 );
	assign w_sys_tmp5694 = (w_sys_tmp5695 < r_run_j_21);
	assign w_sys_tmp5695 = 32'sh00000020;
	assign w_sys_tmp5698 = (w_sys_tmp5699 + r_run_k_20);
	assign w_sys_tmp5699 = (r_run_j_21 * w_sys_tmp5700);
	assign w_sys_tmp5700 = 32'sh00000081;
	assign w_sys_tmp5701 = w_sub00_result_dataout;
	assign w_sys_tmp5702 = (w_sys_tmp5703 + r_run_k_20);
	assign w_sys_tmp5703 = (r_run_copy0_j_131 * w_sys_tmp5700);
	assign w_sys_tmp5705 = (r_run_copy0_j_131 + w_sys_intOne);
	assign w_sys_tmp5706 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp5767 = 32'sh00000021;
	assign w_sys_tmp5768 = ( !w_sys_tmp5769 );
	assign w_sys_tmp5769 = (w_sys_tmp5770 < r_run_j_21);
	assign w_sys_tmp5770 = 32'sh00000040;
	assign w_sys_tmp5772 = (r_run_j_21 - w_sys_tmp5773);
	assign w_sys_tmp5773 = 32'sh0000001f;
	assign w_sys_tmp5775 = (w_sys_tmp5776 + r_run_k_20);
	assign w_sys_tmp5776 = (r_run_copy1_j_133 * w_sys_tmp5777);
	assign w_sys_tmp5777 = 32'sh00000081;
	assign w_sys_tmp5778 = w_sub01_result_dataout;
	assign w_sys_tmp5779 = (w_sys_tmp5780 + r_run_k_20);
	assign w_sys_tmp5780 = (r_run_copy0_j_132 * w_sys_tmp5777);
	assign w_sys_tmp5782 = (r_run_copy0_j_132 + w_sys_intOne);
	assign w_sys_tmp5783 = (r_run_copy1_j_133 + w_sys_intOne);
	assign w_sys_tmp5784 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp5863 = 32'sh00000041;
	assign w_sys_tmp5864 = ( !w_sys_tmp5865 );
	assign w_sys_tmp5865 = (w_sys_tmp5866 < r_run_j_21);
	assign w_sys_tmp5866 = 32'sh00000060;
	assign w_sys_tmp5868 = (r_run_j_21 - w_sys_tmp5869);
	assign w_sys_tmp5869 = 32'sh0000003f;
	assign w_sys_tmp5871 = (w_sys_tmp5872 + r_run_k_20);
	assign w_sys_tmp5872 = (r_run_copy1_j_135 * w_sys_tmp5873);
	assign w_sys_tmp5873 = 32'sh00000081;
	assign w_sys_tmp5874 = w_sub02_result_dataout;
	assign w_sys_tmp5875 = (w_sys_tmp5876 + r_run_k_20);
	assign w_sys_tmp5876 = (r_run_copy0_j_134 * w_sys_tmp5873);
	assign w_sys_tmp5878 = (r_run_copy0_j_134 + w_sys_intOne);
	assign w_sys_tmp5879 = (r_run_copy1_j_135 + w_sys_intOne);
	assign w_sys_tmp5880 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp5959 = 32'sh00000061;
	assign w_sys_tmp5960 = ( !w_sys_tmp5961 );
	assign w_sys_tmp5961 = (w_sys_tmp5962 < r_run_j_21);
	assign w_sys_tmp5962 = 32'sh00000080;
	assign w_sys_tmp5964 = (r_run_j_21 - w_sys_tmp5965);
	assign w_sys_tmp5965 = 32'sh0000005f;
	assign w_sys_tmp5967 = (w_sys_tmp5968 + r_run_k_20);
	assign w_sys_tmp5968 = (r_run_copy1_j_137 * w_sys_tmp5969);
	assign w_sys_tmp5969 = 32'sh00000081;
	assign w_sys_tmp5970 = w_sub03_result_dataout;
	assign w_sys_tmp5971 = (w_sys_tmp5972 + r_run_k_20);
	assign w_sys_tmp5972 = (r_run_copy0_j_136 * w_sys_tmp5969);
	assign w_sys_tmp5974 = (r_run_copy0_j_136 + w_sys_intOne);
	assign w_sys_tmp5975 = (r_run_copy1_j_137 + w_sys_intOne);
	assign w_sys_tmp5976 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6055 = 32'sh00000021;
	assign w_sys_tmp6056 = ( !w_sys_tmp6057 );
	assign w_sys_tmp6057 = (w_sys_tmp6058 < r_run_k_20);
	assign w_sys_tmp6058 = 32'sh00000040;
	assign w_sys_tmp6059 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp6060 = 32'sh00000002;
	assign w_sys_tmp6061 = ( !w_sys_tmp6062 );
	assign w_sys_tmp6062 = (w_sys_tmp6063 < r_run_j_21);
	assign w_sys_tmp6063 = 32'sh00000020;
	assign w_sys_tmp6066 = (w_sys_tmp6067 + r_run_k_20);
	assign w_sys_tmp6067 = (r_run_j_21 * w_sys_tmp6068);
	assign w_sys_tmp6068 = 32'sh00000081;
	assign w_sys_tmp6069 = w_sub04_result_dataout;
	assign w_sys_tmp6070 = (w_sys_tmp6071 + r_run_k_20);
	assign w_sys_tmp6071 = (r_run_copy0_j_138 * w_sys_tmp6068);
	assign w_sys_tmp6073 = (r_run_copy0_j_138 + w_sys_intOne);
	assign w_sys_tmp6074 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6135 = 32'sh00000021;
	assign w_sys_tmp6136 = ( !w_sys_tmp6137 );
	assign w_sys_tmp6137 = (w_sys_tmp6138 < r_run_j_21);
	assign w_sys_tmp6138 = 32'sh00000040;
	assign w_sys_tmp6140 = (r_run_j_21 - w_sys_tmp6141);
	assign w_sys_tmp6141 = 32'sh0000001f;
	assign w_sys_tmp6143 = (w_sys_tmp6144 + r_run_k_20);
	assign w_sys_tmp6144 = (r_run_copy1_j_140 * w_sys_tmp6145);
	assign w_sys_tmp6145 = 32'sh00000081;
	assign w_sys_tmp6146 = w_sub05_result_dataout;
	assign w_sys_tmp6147 = (w_sys_tmp6148 + r_run_k_20);
	assign w_sys_tmp6148 = (r_run_copy0_j_139 * w_sys_tmp6145);
	assign w_sys_tmp6150 = (r_run_copy0_j_139 + w_sys_intOne);
	assign w_sys_tmp6151 = (r_run_copy1_j_140 + w_sys_intOne);
	assign w_sys_tmp6152 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6231 = 32'sh00000041;
	assign w_sys_tmp6232 = ( !w_sys_tmp6233 );
	assign w_sys_tmp6233 = (w_sys_tmp6234 < r_run_j_21);
	assign w_sys_tmp6234 = 32'sh00000060;
	assign w_sys_tmp6236 = (r_run_j_21 - w_sys_tmp6237);
	assign w_sys_tmp6237 = 32'sh0000003f;
	assign w_sys_tmp6239 = (w_sys_tmp6240 + r_run_k_20);
	assign w_sys_tmp6240 = (r_run_copy1_j_142 * w_sys_tmp6241);
	assign w_sys_tmp6241 = 32'sh00000081;
	assign w_sys_tmp6242 = w_sub06_result_dataout;
	assign w_sys_tmp6243 = (w_sys_tmp6244 + r_run_k_20);
	assign w_sys_tmp6244 = (r_run_copy0_j_141 * w_sys_tmp6241);
	assign w_sys_tmp6246 = (r_run_copy0_j_141 + w_sys_intOne);
	assign w_sys_tmp6247 = (r_run_copy1_j_142 + w_sys_intOne);
	assign w_sys_tmp6248 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6327 = 32'sh00000061;
	assign w_sys_tmp6328 = ( !w_sys_tmp6329 );
	assign w_sys_tmp6329 = (w_sys_tmp6330 < r_run_j_21);
	assign w_sys_tmp6330 = 32'sh00000080;
	assign w_sys_tmp6332 = (r_run_j_21 - w_sys_tmp6333);
	assign w_sys_tmp6333 = 32'sh0000005f;
	assign w_sys_tmp6335 = (w_sys_tmp6336 + r_run_k_20);
	assign w_sys_tmp6336 = (r_run_copy1_j_144 * w_sys_tmp6337);
	assign w_sys_tmp6337 = 32'sh00000081;
	assign w_sys_tmp6338 = w_sub07_result_dataout;
	assign w_sys_tmp6339 = (w_sys_tmp6340 + r_run_k_20);
	assign w_sys_tmp6340 = (r_run_copy0_j_143 * w_sys_tmp6337);
	assign w_sys_tmp6342 = (r_run_copy0_j_143 + w_sys_intOne);
	assign w_sys_tmp6343 = (r_run_copy1_j_144 + w_sys_intOne);
	assign w_sys_tmp6344 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6423 = 32'sh00000041;
	assign w_sys_tmp6424 = ( !w_sys_tmp6425 );
	assign w_sys_tmp6425 = (w_sys_tmp6426 < r_run_k_20);
	assign w_sys_tmp6426 = 32'sh00000060;
	assign w_sys_tmp6427 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp6428 = 32'sh00000002;
	assign w_sys_tmp6429 = ( !w_sys_tmp6430 );
	assign w_sys_tmp6430 = (w_sys_tmp6431 < r_run_j_21);
	assign w_sys_tmp6431 = 32'sh00000020;
	assign w_sys_tmp6434 = (w_sys_tmp6435 + r_run_k_20);
	assign w_sys_tmp6435 = (r_run_j_21 * w_sys_tmp6436);
	assign w_sys_tmp6436 = 32'sh00000081;
	assign w_sys_tmp6437 = w_sub08_result_dataout;
	assign w_sys_tmp6438 = (w_sys_tmp6439 + r_run_k_20);
	assign w_sys_tmp6439 = (r_run_copy0_j_145 * w_sys_tmp6436);
	assign w_sys_tmp6441 = (r_run_copy0_j_145 + w_sys_intOne);
	assign w_sys_tmp6442 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6503 = 32'sh00000021;
	assign w_sys_tmp6504 = ( !w_sys_tmp6505 );
	assign w_sys_tmp6505 = (w_sys_tmp6506 < r_run_j_21);
	assign w_sys_tmp6506 = 32'sh00000040;
	assign w_sys_tmp6508 = (r_run_j_21 - w_sys_tmp6509);
	assign w_sys_tmp6509 = 32'sh0000001f;
	assign w_sys_tmp6511 = (w_sys_tmp6512 + r_run_k_20);
	assign w_sys_tmp6512 = (r_run_copy1_j_147 * w_sys_tmp6513);
	assign w_sys_tmp6513 = 32'sh00000081;
	assign w_sys_tmp6514 = w_sub09_result_dataout;
	assign w_sys_tmp6515 = (w_sys_tmp6516 + r_run_k_20);
	assign w_sys_tmp6516 = (r_run_copy0_j_146 * w_sys_tmp6513);
	assign w_sys_tmp6518 = (r_run_copy0_j_146 + w_sys_intOne);
	assign w_sys_tmp6519 = (r_run_copy1_j_147 + w_sys_intOne);
	assign w_sys_tmp6520 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6599 = 32'sh00000041;
	assign w_sys_tmp6600 = ( !w_sys_tmp6601 );
	assign w_sys_tmp6601 = (w_sys_tmp6602 < r_run_j_21);
	assign w_sys_tmp6602 = 32'sh00000060;
	assign w_sys_tmp6604 = (r_run_j_21 - w_sys_tmp6605);
	assign w_sys_tmp6605 = 32'sh0000003f;
	assign w_sys_tmp6607 = (w_sys_tmp6608 + r_run_k_20);
	assign w_sys_tmp6608 = (r_run_copy1_j_149 * w_sys_tmp6609);
	assign w_sys_tmp6609 = 32'sh00000081;
	assign w_sys_tmp6610 = w_sub10_result_dataout;
	assign w_sys_tmp6611 = (w_sys_tmp6612 + r_run_k_20);
	assign w_sys_tmp6612 = (r_run_copy0_j_148 * w_sys_tmp6609);
	assign w_sys_tmp6614 = (r_run_copy0_j_148 + w_sys_intOne);
	assign w_sys_tmp6615 = (r_run_copy1_j_149 + w_sys_intOne);
	assign w_sys_tmp6616 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6695 = 32'sh00000061;
	assign w_sys_tmp6696 = ( !w_sys_tmp6697 );
	assign w_sys_tmp6697 = (w_sys_tmp6698 < r_run_j_21);
	assign w_sys_tmp6698 = 32'sh00000080;
	assign w_sys_tmp6700 = (r_run_j_21 - w_sys_tmp6701);
	assign w_sys_tmp6701 = 32'sh0000005f;
	assign w_sys_tmp6703 = (w_sys_tmp6704 + r_run_k_20);
	assign w_sys_tmp6704 = (r_run_copy1_j_151 * w_sys_tmp6705);
	assign w_sys_tmp6705 = 32'sh00000081;
	assign w_sys_tmp6706 = w_sub11_result_dataout;
	assign w_sys_tmp6707 = (w_sys_tmp6708 + r_run_k_20);
	assign w_sys_tmp6708 = (r_run_copy0_j_150 * w_sys_tmp6705);
	assign w_sys_tmp6710 = (r_run_copy0_j_150 + w_sys_intOne);
	assign w_sys_tmp6711 = (r_run_copy1_j_151 + w_sys_intOne);
	assign w_sys_tmp6712 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6791 = 32'sh00000061;
	assign w_sys_tmp6792 = ( !w_sys_tmp6793 );
	assign w_sys_tmp6793 = (w_sys_tmp6794 < r_run_k_20);
	assign w_sys_tmp6794 = 32'sh00000080;
	assign w_sys_tmp6795 = (r_run_k_20 + w_sys_intOne);
	assign w_sys_tmp6796 = 32'sh00000002;
	assign w_sys_tmp6797 = ( !w_sys_tmp6798 );
	assign w_sys_tmp6798 = (w_sys_tmp6799 < r_run_j_21);
	assign w_sys_tmp6799 = 32'sh00000020;
	assign w_sys_tmp6802 = (w_sys_tmp6803 + r_run_k_20);
	assign w_sys_tmp6803 = (r_run_j_21 * w_sys_tmp6804);
	assign w_sys_tmp6804 = 32'sh00000081;
	assign w_sys_tmp6805 = w_sub12_result_dataout;
	assign w_sys_tmp6806 = (w_sys_tmp6807 + r_run_k_20);
	assign w_sys_tmp6807 = (r_run_copy0_j_152 * w_sys_tmp6804);
	assign w_sys_tmp6809 = (r_run_copy0_j_152 + w_sys_intOne);
	assign w_sys_tmp6810 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6871 = 32'sh00000021;
	assign w_sys_tmp6872 = ( !w_sys_tmp6873 );
	assign w_sys_tmp6873 = (w_sys_tmp6874 < r_run_j_21);
	assign w_sys_tmp6874 = 32'sh00000040;
	assign w_sys_tmp6876 = (r_run_j_21 - w_sys_tmp6877);
	assign w_sys_tmp6877 = 32'sh0000001f;
	assign w_sys_tmp6879 = (w_sys_tmp6880 + r_run_k_20);
	assign w_sys_tmp6880 = (r_run_copy1_j_154 * w_sys_tmp6881);
	assign w_sys_tmp6881 = 32'sh00000081;
	assign w_sys_tmp6882 = w_sub13_result_dataout;
	assign w_sys_tmp6883 = (w_sys_tmp6884 + r_run_k_20);
	assign w_sys_tmp6884 = (r_run_copy0_j_153 * w_sys_tmp6881);
	assign w_sys_tmp6886 = (r_run_copy0_j_153 + w_sys_intOne);
	assign w_sys_tmp6887 = (r_run_copy1_j_154 + w_sys_intOne);
	assign w_sys_tmp6888 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp6967 = 32'sh00000041;
	assign w_sys_tmp6968 = ( !w_sys_tmp6969 );
	assign w_sys_tmp6969 = (w_sys_tmp6970 < r_run_j_21);
	assign w_sys_tmp6970 = 32'sh00000060;
	assign w_sys_tmp6972 = (r_run_j_21 - w_sys_tmp6973);
	assign w_sys_tmp6973 = 32'sh0000003f;
	assign w_sys_tmp6975 = (w_sys_tmp6976 + r_run_k_20);
	assign w_sys_tmp6976 = (r_run_copy1_j_156 * w_sys_tmp6977);
	assign w_sys_tmp6977 = 32'sh00000081;
	assign w_sys_tmp6978 = w_sub14_result_dataout;
	assign w_sys_tmp6979 = (w_sys_tmp6980 + r_run_k_20);
	assign w_sys_tmp6980 = (r_run_copy0_j_155 * w_sys_tmp6977);
	assign w_sys_tmp6982 = (r_run_copy0_j_155 + w_sys_intOne);
	assign w_sys_tmp6983 = (r_run_copy1_j_156 + w_sys_intOne);
	assign w_sys_tmp6984 = (r_run_j_21 + w_sys_intOne);
	assign w_sys_tmp7063 = 32'sh00000061;
	assign w_sys_tmp7064 = ( !w_sys_tmp7065 );
	assign w_sys_tmp7065 = (w_sys_tmp7066 < r_run_j_21);
	assign w_sys_tmp7066 = 32'sh00000080;
	assign w_sys_tmp7068 = (r_run_j_21 - w_sys_tmp7069);
	assign w_sys_tmp7069 = 32'sh0000005f;
	assign w_sys_tmp7071 = (w_sys_tmp7072 + r_run_k_20);
	assign w_sys_tmp7072 = (r_run_copy1_j_158 * w_sys_tmp7073);
	assign w_sys_tmp7073 = 32'sh00000081;
	assign w_sys_tmp7074 = w_sub15_result_dataout;
	assign w_sys_tmp7075 = (w_sys_tmp7076 + r_run_k_20);
	assign w_sys_tmp7076 = (r_run_copy0_j_157 * w_sys_tmp7073);
	assign w_sys_tmp7078 = (r_run_copy0_j_157 + w_sys_intOne);
	assign w_sys_tmp7079 = (r_run_copy1_j_158 + w_sys_intOne);
	assign w_sys_tmp7080 = (r_run_j_21 + w_sys_intOne);


	sub09
		sub09_inst(
			.i_fld_T_0_addr_0 (w_sub09_T_addr),
			.i_fld_T_0_datain_0 (w_sub09_T_datain),
			.o_fld_T_0_dataout_0 (w_sub09_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub09_T_r_w),
			.i_fld_U_2_addr_0 (w_sub09_U_addr),
			.i_fld_U_2_datain_0 (w_sub09_U_datain),
			.o_fld_U_2_dataout_0 (w_sub09_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub09_U_r_w),
			.i_fld_V_1_addr_0 (w_sub09_V_addr),
			.i_fld_V_1_datain_0 (w_sub09_V_datain),
			.o_fld_V_1_dataout_0 (w_sub09_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub09_V_r_w),
			.i_fld_result_3_addr_0 (w_sub09_result_addr),
			.i_fld_result_3_datain_0 (w_sub09_result_datain),
			.o_fld_result_3_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub09_result_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_T_0_addr_0 (w_sub08_T_addr),
			.i_fld_T_0_datain_0 (w_sub08_T_datain),
			.o_fld_T_0_dataout_0 (w_sub08_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub08_T_r_w),
			.i_fld_U_2_addr_0 (w_sub08_U_addr),
			.i_fld_U_2_datain_0 (w_sub08_U_datain),
			.o_fld_U_2_dataout_0 (w_sub08_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub08_U_r_w),
			.i_fld_V_1_addr_0 (w_sub08_V_addr),
			.i_fld_V_1_datain_0 (w_sub08_V_datain),
			.o_fld_V_1_dataout_0 (w_sub08_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub08_V_r_w),
			.i_fld_result_3_addr_0 (w_sub08_result_addr),
			.i_fld_result_3_datain_0 (w_sub08_result_datain),
			.o_fld_result_3_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub08_result_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_T_0_addr_0 (w_sub12_T_addr),
			.i_fld_T_0_datain_0 (w_sub12_T_datain),
			.o_fld_T_0_dataout_0 (w_sub12_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub12_T_r_w),
			.i_fld_U_2_addr_0 (w_sub12_U_addr),
			.i_fld_U_2_datain_0 (w_sub12_U_datain),
			.o_fld_U_2_dataout_0 (w_sub12_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub12_U_r_w),
			.i_fld_V_1_addr_0 (w_sub12_V_addr),
			.i_fld_V_1_datain_0 (w_sub12_V_datain),
			.o_fld_V_1_dataout_0 (w_sub12_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub12_V_r_w),
			.i_fld_result_3_addr_0 (w_sub12_result_addr),
			.i_fld_result_3_datain_0 (w_sub12_result_datain),
			.o_fld_result_3_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub12_result_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_T_0_addr_0 (w_sub03_T_addr),
			.i_fld_T_0_datain_0 (w_sub03_T_datain),
			.o_fld_T_0_dataout_0 (w_sub03_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub03_T_r_w),
			.i_fld_U_2_addr_0 (w_sub03_U_addr),
			.i_fld_U_2_datain_0 (w_sub03_U_datain),
			.o_fld_U_2_dataout_0 (w_sub03_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub03_U_r_w),
			.i_fld_V_1_addr_0 (w_sub03_V_addr),
			.i_fld_V_1_datain_0 (w_sub03_V_datain),
			.o_fld_V_1_dataout_0 (w_sub03_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub03_V_r_w),
			.i_fld_result_3_addr_0 (w_sub03_result_addr),
			.i_fld_result_3_datain_0 (w_sub03_result_datain),
			.o_fld_result_3_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub03_result_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_T_0_addr_0 (w_sub02_T_addr),
			.i_fld_T_0_datain_0 (w_sub02_T_datain),
			.o_fld_T_0_dataout_0 (w_sub02_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub02_T_r_w),
			.i_fld_U_2_addr_0 (w_sub02_U_addr),
			.i_fld_U_2_datain_0 (w_sub02_U_datain),
			.o_fld_U_2_dataout_0 (w_sub02_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub02_U_r_w),
			.i_fld_V_1_addr_0 (w_sub02_V_addr),
			.i_fld_V_1_datain_0 (w_sub02_V_datain),
			.o_fld_V_1_dataout_0 (w_sub02_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub02_V_r_w),
			.i_fld_result_3_addr_0 (w_sub02_result_addr),
			.i_fld_result_3_datain_0 (w_sub02_result_datain),
			.o_fld_result_3_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub02_result_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_T_0_addr_0 (w_sub11_T_addr),
			.i_fld_T_0_datain_0 (w_sub11_T_datain),
			.o_fld_T_0_dataout_0 (w_sub11_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub11_T_r_w),
			.i_fld_U_2_addr_0 (w_sub11_U_addr),
			.i_fld_U_2_datain_0 (w_sub11_U_datain),
			.o_fld_U_2_dataout_0 (w_sub11_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub11_U_r_w),
			.i_fld_V_1_addr_0 (w_sub11_V_addr),
			.i_fld_V_1_datain_0 (w_sub11_V_datain),
			.o_fld_V_1_dataout_0 (w_sub11_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub11_V_r_w),
			.i_fld_result_3_addr_0 (w_sub11_result_addr),
			.i_fld_result_3_datain_0 (w_sub11_result_datain),
			.o_fld_result_3_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub11_result_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_T_0_addr_0 (w_sub14_T_addr),
			.i_fld_T_0_datain_0 (w_sub14_T_datain),
			.o_fld_T_0_dataout_0 (w_sub14_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub14_T_r_w),
			.i_fld_U_2_addr_0 (w_sub14_U_addr),
			.i_fld_U_2_datain_0 (w_sub14_U_datain),
			.o_fld_U_2_dataout_0 (w_sub14_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub14_U_r_w),
			.i_fld_V_1_addr_0 (w_sub14_V_addr),
			.i_fld_V_1_datain_0 (w_sub14_V_datain),
			.o_fld_V_1_dataout_0 (w_sub14_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub14_V_r_w),
			.i_fld_result_3_addr_0 (w_sub14_result_addr),
			.i_fld_result_3_datain_0 (w_sub14_result_datain),
			.o_fld_result_3_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub14_result_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_T_0_addr_0 (w_sub01_T_addr),
			.i_fld_T_0_datain_0 (w_sub01_T_datain),
			.o_fld_T_0_dataout_0 (w_sub01_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub01_T_r_w),
			.i_fld_U_2_addr_0 (w_sub01_U_addr),
			.i_fld_U_2_datain_0 (w_sub01_U_datain),
			.o_fld_U_2_dataout_0 (w_sub01_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub01_U_r_w),
			.i_fld_V_1_addr_0 (w_sub01_V_addr),
			.i_fld_V_1_datain_0 (w_sub01_V_datain),
			.o_fld_V_1_dataout_0 (w_sub01_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub01_V_r_w),
			.i_fld_result_3_addr_0 (w_sub01_result_addr),
			.i_fld_result_3_datain_0 (w_sub01_result_datain),
			.o_fld_result_3_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub01_result_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_T_0_addr_0 (w_sub13_T_addr),
			.i_fld_T_0_datain_0 (w_sub13_T_datain),
			.o_fld_T_0_dataout_0 (w_sub13_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub13_T_r_w),
			.i_fld_U_2_addr_0 (w_sub13_U_addr),
			.i_fld_U_2_datain_0 (w_sub13_U_datain),
			.o_fld_U_2_dataout_0 (w_sub13_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub13_U_r_w),
			.i_fld_V_1_addr_0 (w_sub13_V_addr),
			.i_fld_V_1_datain_0 (w_sub13_V_datain),
			.o_fld_V_1_dataout_0 (w_sub13_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub13_V_r_w),
			.i_fld_result_3_addr_0 (w_sub13_result_addr),
			.i_fld_result_3_datain_0 (w_sub13_result_datain),
			.o_fld_result_3_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub13_result_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_T_0_addr_0 (w_sub00_T_addr),
			.i_fld_T_0_datain_0 (w_sub00_T_datain),
			.o_fld_T_0_dataout_0 (w_sub00_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub00_T_r_w),
			.i_fld_U_2_addr_0 (w_sub00_U_addr),
			.i_fld_U_2_datain_0 (w_sub00_U_datain),
			.o_fld_U_2_dataout_0 (w_sub00_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub00_U_r_w),
			.i_fld_V_1_addr_0 (w_sub00_V_addr),
			.i_fld_V_1_datain_0 (w_sub00_V_datain),
			.o_fld_V_1_dataout_0 (w_sub00_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub00_V_r_w),
			.i_fld_result_3_addr_0 (w_sub00_result_addr),
			.i_fld_result_3_datain_0 (w_sub00_result_datain),
			.o_fld_result_3_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub00_result_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_T_0_addr_0 (w_sub07_T_addr),
			.i_fld_T_0_datain_0 (w_sub07_T_datain),
			.o_fld_T_0_dataout_0 (w_sub07_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub07_T_r_w),
			.i_fld_U_2_addr_0 (w_sub07_U_addr),
			.i_fld_U_2_datain_0 (w_sub07_U_datain),
			.o_fld_U_2_dataout_0 (w_sub07_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub07_U_r_w),
			.i_fld_V_1_addr_0 (w_sub07_V_addr),
			.i_fld_V_1_datain_0 (w_sub07_V_datain),
			.o_fld_V_1_dataout_0 (w_sub07_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub07_V_r_w),
			.i_fld_result_3_addr_0 (w_sub07_result_addr),
			.i_fld_result_3_datain_0 (w_sub07_result_datain),
			.o_fld_result_3_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub07_result_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_T_0_addr_0 (w_sub06_T_addr),
			.i_fld_T_0_datain_0 (w_sub06_T_datain),
			.o_fld_T_0_dataout_0 (w_sub06_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub06_T_r_w),
			.i_fld_U_2_addr_0 (w_sub06_U_addr),
			.i_fld_U_2_datain_0 (w_sub06_U_datain),
			.o_fld_U_2_dataout_0 (w_sub06_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub06_U_r_w),
			.i_fld_V_1_addr_0 (w_sub06_V_addr),
			.i_fld_V_1_datain_0 (w_sub06_V_datain),
			.o_fld_V_1_dataout_0 (w_sub06_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub06_V_r_w),
			.i_fld_result_3_addr_0 (w_sub06_result_addr),
			.i_fld_result_3_datain_0 (w_sub06_result_datain),
			.o_fld_result_3_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub06_result_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_T_0_addr_0 (w_sub15_T_addr),
			.i_fld_T_0_datain_0 (w_sub15_T_datain),
			.o_fld_T_0_dataout_0 (w_sub15_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub15_T_r_w),
			.i_fld_U_2_addr_0 (w_sub15_U_addr),
			.i_fld_U_2_datain_0 (w_sub15_U_datain),
			.o_fld_U_2_dataout_0 (w_sub15_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub15_U_r_w),
			.i_fld_V_1_addr_0 (w_sub15_V_addr),
			.i_fld_V_1_datain_0 (w_sub15_V_datain),
			.o_fld_V_1_dataout_0 (w_sub15_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub15_V_r_w),
			.i_fld_result_3_addr_0 (w_sub15_result_addr),
			.i_fld_result_3_datain_0 (w_sub15_result_datain),
			.o_fld_result_3_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub15_result_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_T_0_addr_0 (w_sub05_T_addr),
			.i_fld_T_0_datain_0 (w_sub05_T_datain),
			.o_fld_T_0_dataout_0 (w_sub05_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub05_T_r_w),
			.i_fld_U_2_addr_0 (w_sub05_U_addr),
			.i_fld_U_2_datain_0 (w_sub05_U_datain),
			.o_fld_U_2_dataout_0 (w_sub05_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub05_U_r_w),
			.i_fld_V_1_addr_0 (w_sub05_V_addr),
			.i_fld_V_1_datain_0 (w_sub05_V_datain),
			.o_fld_V_1_dataout_0 (w_sub05_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub05_V_r_w),
			.i_fld_result_3_addr_0 (w_sub05_result_addr),
			.i_fld_result_3_datain_0 (w_sub05_result_datain),
			.o_fld_result_3_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub05_result_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_T_0_addr_0 (w_sub04_T_addr),
			.i_fld_T_0_datain_0 (w_sub04_T_datain),
			.o_fld_T_0_dataout_0 (w_sub04_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub04_T_r_w),
			.i_fld_U_2_addr_0 (w_sub04_U_addr),
			.i_fld_U_2_datain_0 (w_sub04_U_datain),
			.o_fld_U_2_dataout_0 (w_sub04_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub04_U_r_w),
			.i_fld_V_1_addr_0 (w_sub04_V_addr),
			.i_fld_V_1_datain_0 (w_sub04_V_datain),
			.o_fld_V_1_dataout_0 (w_sub04_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub04_V_r_w),
			.i_fld_result_3_addr_0 (w_sub04_result_addr),
			.i_fld_result_3_datain_0 (w_sub04_result_datain),
			.o_fld_result_3_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub04_result_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_T_0_addr_0 (w_sub10_T_addr),
			.i_fld_T_0_datain_0 (w_sub10_T_datain),
			.o_fld_T_0_dataout_0 (w_sub10_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub10_T_r_w),
			.i_fld_U_2_addr_0 (w_sub10_U_addr),
			.i_fld_U_2_datain_0 (w_sub10_U_datain),
			.o_fld_U_2_dataout_0 (w_sub10_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub10_U_r_w),
			.i_fld_V_1_addr_0 (w_sub10_V_addr),
			.i_fld_V_1_datain_0 (w_sub10_V_datain),
			.o_fld_V_1_dataout_0 (w_sub10_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub10_V_r_w),
			.i_fld_result_3_addr_0 (w_sub10_result_addr),
			.i_fld_result_3_datain_0 (w_sub10_result_datain),
			.o_fld_result_3_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub10_result_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_V_3(
			.clk (clock),
			.ce_0 (w_fld_V_3_ce_0),
			.addr_0 (w_fld_V_3_addr_0),
			.datain_0 (w_fld_V_3_datain_0),
			.dataout_0 (w_fld_V_3_dataout_0),
			.r_w_0 (w_fld_V_3_r_w_0),
			.ce_1 (w_fld_V_3_ce_1),
			.addr_1 (r_fld_V_3_addr_1),
			.datain_1 (r_fld_V_3_datain_1),
			.dataout_1 (w_fld_V_3_dataout_1),
			.r_w_1 (r_fld_V_3_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp39;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp129[31], w_sys_tmp129[30:0] };

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp129[31], w_sys_tmp129[30:0] };

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h7<=r_sys_run_step && r_sys_run_step<=7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'hf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_27;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h16)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp37;

									end
									else
									if((r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h16)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_32;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp38;

									end
									else
									if((r_sys_run_step==7'h15) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((7'h7<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp20;

									end
									else
									if((r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp21;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						9'h12f: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 9'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h0: begin
							r_sys_run_phase <= 9'h2;
						end

						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h4;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h5;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13) ? 9'h9 : 9'hf);

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h5;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'ha;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp16) ? 9'hd : 9'h6);

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h20)) begin
										r_sys_run_phase <= 9'ha;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h10;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp227) ? 9'h14 : 9'h2c);

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h10;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h15;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp231) ? 9'h18 : 9'h1a);

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h15;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h1b;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp446) ? 9'h1e : 9'h20);

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h1b;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h21;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp661) ? 9'h24 : 9'h26);

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h21;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h27;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp876) ? 9'h2a : 9'h11);

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h27;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h2d;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1091) ? 9'h31 : 9'h49);

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h2d;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h32;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1095) ? 9'h35 : 9'h37);

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h32;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h38;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1310) ? 9'h3b : 9'h3d);

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h38;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h3e;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1525) ? 9'h41 : 9'h43);

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h3e;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h44;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1740) ? 9'h47 : 9'h2e);

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h44;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h4a;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1955) ? 9'h4e : 9'h66);

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h4a;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h4f;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1959) ? 9'h52 : 9'h54);

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h4f;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h55;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2174) ? 9'h58 : 9'h5a);

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h55;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h5b;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2389) ? 9'h5e : 9'h60);

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h5b;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h61;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2604) ? 9'h64 : 9'h4b);

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h61;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h67;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2819) ? 9'h6b : 9'h83);

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h67;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h6c;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2823) ? 9'h6f : 9'h71);

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h6c;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h72;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3038) ? 9'h75 : 9'h77);

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h72;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h78;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3253) ? 9'h7b : 9'h7d);

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h78;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h7e;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3468) ? 9'h81 : 9'h68);

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h7e;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h84;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3682) ? 9'h87 : 9'hbb);

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h84;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 9'h89;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 9'h8b;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h8c;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3686) ? 9'h8f : 9'h91);

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_phase <= 9'h8c;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h92;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3726) ? 9'h95 : 9'h97);

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_phase <= 9'h92;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h98;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3766) ? 9'h9b : 9'h9d);

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_phase <= 9'h98;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h9e;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3806) ? 9'ha1 : 9'ha3);

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_phase <= 9'h9e;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'ha4;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3846) ? 9'ha7 : 9'ha9);

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3d)) begin
										r_sys_run_phase <= 9'ha4;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'haa;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4347) ? 9'had : 9'haf);

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_phase <= 9'haa;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hb0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4794) ? 9'hb3 : 9'hb5);

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_phase <= 9'hb0;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hb6;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5241) ? 9'hb9 : 9'h85);

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_phase <= 9'hb6;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hbc;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5688) ? 9'hc0 : 9'hd8);

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hbc;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hc1;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5693) ? 9'hc4 : 9'hc6);

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hc1;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hc7;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5768) ? 9'hca : 9'hcc);

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hc7;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hcd;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5864) ? 9'hd0 : 9'hd2);

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hcd;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hd3;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5960) ? 9'hd6 : 9'hbd);

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hd3;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hd9;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6056) ? 9'hdd : 9'hf5);

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hd9;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hde;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6061) ? 9'he1 : 9'he3);

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hde;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'he4;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6136) ? 9'he7 : 9'he9);

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'he4;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hea;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6232) ? 9'hed : 9'hef);

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hea;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hf0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6328) ? 9'hf3 : 9'hda);

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hf0;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hf6;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6424) ? 9'hfa : 9'h112);

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hf6;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'hfb;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6429) ? 9'hfe : 9'h100);

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'hfb;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h101;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6504) ? 9'h104 : 9'h106);

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h101;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h107;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6600) ? 9'h10a : 9'h10c);

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h107;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h10d;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6696) ? 9'h110 : 9'hf7);

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h10d;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h113;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6792) ? 9'h117 : 9'h12f);

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h113;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h118;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6797) ? 9'h11b : 9'h11d);

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h118;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h11e;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6872) ? 9'h121 : 9'h123);

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h11e;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h124;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6968) ? 9'h127 : 9'h129);

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h124;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 9'h12a;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7064) ? 9'h12d : 9'h114);

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_phase <= 9'h12a;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sys_run_phase <= 9'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h20)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h20)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h6c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h72: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h78: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h89: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h8c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h92: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h98: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h9e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'ha4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3d)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'haa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hb6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5b)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hbc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hc1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hc7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hcd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hd9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hf0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hf6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h118: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h11e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h124: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h12a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						9'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						9'h12f: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp23[14:0] );

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp256[14:0] );

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp471[14:0] );

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp686[14:0] );

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp901[14:0] );

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1120[14:0] );

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1335[14:0] );

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1550[14:0] );

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1765[14:0] );

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1984[14:0] );

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2199[14:0] );

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2414[14:0] );

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2629[14:0] );

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2848[14:0] );

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3063[14:0] );

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3278[14:0] );

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3493[14:0] );

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp5698[14:0] );

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp5775[14:0] );

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp5871[14:0] );

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp5967[14:0] );

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6066[14:0] );

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6143[14:0] );

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6239[14:0] );

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6335[14:0] );

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6434[14:0] );

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6511[14:0] );

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6607[14:0] );

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6703[14:0] );

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6802[14:0] );

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6879[14:0] );

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6975[14:0] );

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7071[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp5701;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp5778;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp5874;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp5970;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6069;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6146;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6242;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6338;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6437;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6514;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6610;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6706;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6805;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6882;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp6978;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp7074;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12f: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp28[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h12f: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp33[14:0] );

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp240[14:0] );

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp455[14:0] );

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp670[14:0] );

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp885[14:0] );

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1104[14:0] );

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1319[14:0] );

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1534[14:0] );

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1749[14:0] );

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1968[14:0] );

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2183[14:0] );

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2398[14:0] );

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2613[14:0] );

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2832[14:0] );

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3047[14:0] );

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3262[14:0] );

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3477[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp19;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp42[14:0] );

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp248[14:0] );

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp463[14:0] );

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp678[14:0] );

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp893[14:0] );

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1112[14:0] );

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1327[14:0] );

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1542[14:0] );

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1757[14:0] );

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1976[14:0] );

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2191[14:0] );

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2406[14:0] );

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2621[14:0] );

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2840[14:0] );

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3055[14:0] );

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3270[14:0] );

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3485[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_fld_V_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp15;

									end
								end

							endcase
						end

						9'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp230;

									end
								end

							endcase
						end

						9'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp1090;

									end
								end

							endcase
						end

						9'h2e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp1094;

									end
								end

							endcase
						end

						9'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp1954;

									end
								end

							endcase
						end

						9'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp1958;

									end
								end

							endcase
						end

						9'h66: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp2818;

									end
								end

							endcase
						end

						9'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp2822;

									end
								end

							endcase
						end

						9'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp3685;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_run_k_20 <= w_sys_tmp3724;

									end
								end

							endcase
						end

						9'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp3725;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_run_k_20 <= w_sys_tmp3764;

									end
								end

							endcase
						end

						9'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp3765;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_run_k_20 <= w_sys_tmp3804;

									end
								end

							endcase
						end

						9'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp3805;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_run_k_20 <= w_sys_tmp3844;

									end
								end

							endcase
						end

						9'hbb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp5687;

									end
								end

							endcase
						end

						9'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp5691;

									end
								end

							endcase
						end

						9'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp6055;

									end
								end

							endcase
						end

						9'hda: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp6059;

									end
								end

							endcase
						end

						9'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp6423;

									end
								end

							endcase
						end

						9'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp6427;

									end
								end

							endcase
						end

						9'h112: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp6791;

									end
								end

							endcase
						end

						9'h114: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_20 <= w_sys_tmp6795;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp49;

									end
								end

							endcase
						end

						9'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp264;

									end
								end

							endcase
						end

						9'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp445;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp479;

									end
								end

							endcase
						end

						9'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp660;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp694;

									end
								end

							endcase
						end

						9'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp875;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp909;

									end
								end

							endcase
						end

						9'h31: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp1128;

									end
								end

							endcase
						end

						9'h37: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp1309;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp1343;

									end
								end

							endcase
						end

						9'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp1524;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp1558;

									end
								end

							endcase
						end

						9'h43: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp1739;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp1773;

									end
								end

							endcase
						end

						9'h4e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp1992;

									end
								end

							endcase
						end

						9'h54: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp2173;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp2207;

									end
								end

							endcase
						end

						9'h5a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp2388;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp2422;

									end
								end

							endcase
						end

						9'h60: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp2603;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp2637;

									end
								end

							endcase
						end

						9'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp2856;

									end
								end

							endcase
						end

						9'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp3037;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp3071;

									end
								end

							endcase
						end

						9'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp3252;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp3286;

									end
								end

							endcase
						end

						9'h7d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp3467;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp3501;

									end
								end

							endcase
						end

						9'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp3845;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32)) begin
										r_run_j_21 <= w_sys_tmp3919;

									end
								end

							endcase
						end

						9'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp4346;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_j_21 <= w_sys_tmp4414;

									end
								end

							endcase
						end

						9'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp4793;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_j_21 <= w_sys_tmp4861;

									end
								end

							endcase
						end

						9'hb5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp5240;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_j_21 <= w_sys_tmp5308;

									end
								end

							endcase
						end

						9'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp5692;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp5706;

									end
								end

							endcase
						end

						9'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp5767;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp5784;

									end
								end

							endcase
						end

						9'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp5863;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp5880;

									end
								end

							endcase
						end

						9'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp5959;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp5976;

									end
								end

							endcase
						end

						9'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6060;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp6074;

									end
								end

							endcase
						end

						9'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6135;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp6152;

									end
								end

							endcase
						end

						9'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6231;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp6248;

									end
								end

							endcase
						end

						9'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6327;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp6344;

									end
								end

							endcase
						end

						9'hfa: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6428;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp6442;

									end
								end

							endcase
						end

						9'h100: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6503;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp6520;

									end
								end

							endcase
						end

						9'h106: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6599;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp6616;

									end
								end

							endcase
						end

						9'h10c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6695;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp6712;

									end
								end

							endcase
						end

						9'h117: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6796;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_j_21 <= w_sys_tmp6810;

									end
								end

							endcase
						end

						9'h11d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6871;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp6888;

									end
								end

							endcase
						end

						9'h123: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp6967;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp6984;

									end
								end

							endcase
						end

						9'h129: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_21 <= w_sys_tmp7063;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_21 <= w_sys_tmp7080;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h83: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_22 <= w_sys_intOne;

									end
								end

							endcase
						end

						9'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_22 <= w_sys_tmp3684;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_mx_23 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_my_24 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dt_25 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dx_26 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dy_27 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r1_28 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r2_29 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r3_30 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r4_31 <= w_sys_tmp12;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14)) begin
										r_run_YY_32 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h11)) begin
										r_run_YY_32 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_kx_33 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_ky_34 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_nlast_35 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_tmpj_36 <= w_sys_tmp4351;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_tmpj_36 <= w_sys_tmp4798;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_run_tmpj_36 <= w_sys_tmp5245;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp5772;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp5868;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp5964;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp6140;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp6236;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp6332;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp6508;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp6604;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp6700;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp6876;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp6972;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_tmpj_36 <= w_sys_tmp7068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_37 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_37 <= w_sys_tmp46;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_38 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_run_copy1_j_38 <= w_sys_tmp47;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_39 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_39 <= w_sys_tmp48;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_40 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_40 <= w_sys_tmp259;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_41 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_41 <= w_sys_tmp260;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_42 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_42 <= w_sys_tmp261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_43 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_43 <= w_sys_tmp262;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_44 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_44 <= w_sys_tmp263;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_45 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_45 <= w_sys_tmp474;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_46 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_46 <= w_sys_tmp475;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_47 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_47 <= w_sys_tmp476;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_48 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_48 <= w_sys_tmp477;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_49 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_49 <= w_sys_tmp478;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_50 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_50 <= w_sys_tmp689;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_51 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_51 <= w_sys_tmp690;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_52 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_52 <= w_sys_tmp691;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_53 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_53 <= w_sys_tmp692;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_54 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_54 <= w_sys_tmp693;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_55 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_55 <= w_sys_tmp904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_56 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_56 <= w_sys_tmp905;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_57 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_57 <= w_sys_tmp906;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_58 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_58 <= w_sys_tmp907;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_59 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_59 <= w_sys_tmp908;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_60 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_60 <= w_sys_tmp1123;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_61 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_61 <= w_sys_tmp1124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_62 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_62 <= w_sys_tmp1125;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_63 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_63 <= w_sys_tmp1126;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h31: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_64 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_64 <= w_sys_tmp1127;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_65 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_65 <= w_sys_tmp1338;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_66 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_66 <= w_sys_tmp1339;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_67 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_67 <= w_sys_tmp1340;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_68 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_68 <= w_sys_tmp1341;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h37: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_69 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_69 <= w_sys_tmp1342;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_70 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_70 <= w_sys_tmp1553;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_71 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_71 <= w_sys_tmp1554;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_72 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_72 <= w_sys_tmp1555;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_73 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_73 <= w_sys_tmp1556;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_74 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_74 <= w_sys_tmp1557;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_75 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_75 <= w_sys_tmp1768;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_76 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_76 <= w_sys_tmp1769;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_77 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_77 <= w_sys_tmp1770;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_78 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_78 <= w_sys_tmp1771;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h43: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_79 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_79 <= w_sys_tmp1772;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_80 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_80 <= w_sys_tmp1987;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_81 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_81 <= w_sys_tmp1988;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_82 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_82 <= w_sys_tmp1989;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_83 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_83 <= w_sys_tmp1990;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h4e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_84 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_84 <= w_sys_tmp1991;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_85 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_85 <= w_sys_tmp2202;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_86 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_86 <= w_sys_tmp2203;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_87 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_87 <= w_sys_tmp2204;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_88 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_88 <= w_sys_tmp2205;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h54: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_89 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_89 <= w_sys_tmp2206;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_90 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_90 <= w_sys_tmp2417;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_91 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_91 <= w_sys_tmp2418;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_92 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_92 <= w_sys_tmp2419;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_93 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_93 <= w_sys_tmp2420;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_94 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_94 <= w_sys_tmp2421;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_95 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_95 <= w_sys_tmp2632;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_96 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_96 <= w_sys_tmp2633;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_97 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_97 <= w_sys_tmp2634;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_98 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_98 <= w_sys_tmp2635;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h60: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_99 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_99 <= w_sys_tmp2636;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_100 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_100 <= w_sys_tmp2851;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_101 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_101 <= w_sys_tmp2852;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_102 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_102 <= w_sys_tmp2853;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_103 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_103 <= w_sys_tmp2854;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_104 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_104 <= w_sys_tmp2855;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_105 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_105 <= w_sys_tmp3066;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_106 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_106 <= w_sys_tmp3067;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_107 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_107 <= w_sys_tmp3068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_108 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_108 <= w_sys_tmp3069;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h71: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_109 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_109 <= w_sys_tmp3070;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_110 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_110 <= w_sys_tmp3281;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_111 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_111 <= w_sys_tmp3282;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_112 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_112 <= w_sys_tmp3283;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_113 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_113 <= w_sys_tmp3284;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h77: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_114 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_114 <= w_sys_tmp3285;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_115 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_115 <= w_sys_tmp3496;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_116 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_116 <= w_sys_tmp3497;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_117 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_117 <= w_sys_tmp3498;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_118 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy3_j_118 <= w_sys_tmp3499;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_119 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy4_j_119 <= w_sys_tmp3500;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_120 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h3b)) begin
										r_run_copy0_j_120 <= w_sys_tmp3908;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_121 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h3d)) begin
										r_run_copy1_j_121 <= w_sys_tmp3909;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_122 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_run_copy2_j_122 <= w_sys_tmp3910;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_123 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3a)) begin
										r_run_copy3_j_123 <= w_sys_tmp3911;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_124 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h37)) begin
										r_run_copy4_j_124 <= w_sys_tmp3912;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy5_j_125 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h39)) begin
										r_run_copy5_j_125 <= w_sys_tmp3913;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy6_j_126 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h34)) begin
										r_run_copy6_j_126 <= w_sys_tmp3914;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy7_j_127 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_run_copy7_j_127 <= w_sys_tmp3915;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy8_j_128 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33)) begin
										r_run_copy8_j_128 <= w_sys_tmp3916;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy9_j_129 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35)) begin
										r_run_copy9_j_129 <= w_sys_tmp3917;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy10_j_130 <= r_run_j_21;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h30)) begin
										r_run_copy10_j_130 <= w_sys_tmp3918;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_131 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_131 <= w_sys_tmp5705;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_132 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_132 <= w_sys_tmp5782;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hc6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_133 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_133 <= w_sys_tmp5783;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hcc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_134 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_134 <= w_sys_tmp5878;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hcc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_135 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_135 <= w_sys_tmp5879;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_136 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_136 <= w_sys_tmp5974;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_137 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_137 <= w_sys_tmp5975;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_138 <= r_run_j_21;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_138 <= w_sys_tmp6073;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_139 <= r_run_j_21;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_139 <= w_sys_tmp6150;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_140 <= r_run_j_21;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_140 <= w_sys_tmp6151;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_141 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_141 <= w_sys_tmp6246;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'he9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_142 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_142 <= w_sys_tmp6247;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_143 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_143 <= w_sys_tmp6342;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_144 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_144 <= w_sys_tmp6343;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hfa: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_145 <= r_run_j_21;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_145 <= w_sys_tmp6441;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h100: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_146 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_146 <= w_sys_tmp6518;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h100: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_147 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_147 <= w_sys_tmp6519;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h106: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_148 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_148 <= w_sys_tmp6614;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h106: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_149 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_149 <= w_sys_tmp6615;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h10c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_150 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_150 <= w_sys_tmp6710;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h10c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_151 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_151 <= w_sys_tmp6711;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h117: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_152 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_152 <= w_sys_tmp6809;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h11d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_153 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_153 <= w_sys_tmp6886;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h11d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_154 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_154 <= w_sys_tmp6887;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h123: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_155 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_155 <= w_sys_tmp6982;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h123: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_156 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_156 <= w_sys_tmp6983;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h129: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_157 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_157 <= w_sys_tmp7078;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h129: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_158 <= r_run_j_21;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_run_copy1_j_158 <= w_sys_tmp7079;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp2195[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_T_datain <= w_sys_tmp2198;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp2187[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_V_datain <= w_sys_tmp2190;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp2179[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_U_datain <= w_sys_tmp2182;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h58: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub09_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3783[14:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3777[14:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3771[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3774[14:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4395[14:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h59)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4405[14:0] );

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4385[14:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp4379[14:0] );

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp6515[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub09_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub09_result_datain <= w_sys_tmp3779;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub09_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub09_result_datain <= w_sys_tmp4358;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h57) || (r_sys_run_step==7'h58)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h59)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp1980[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_T_datain <= w_sys_tmp1983;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1972[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_V_datain <= w_sys_tmp1975;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1964[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_U_datain <= w_sys_tmp1967;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h52: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3780[14:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3771[14:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3a)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3890[14:0] );

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h39)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3880[14:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h34)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3875[14:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h3b)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3904[14:0] );

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp6438[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_datain <= w_sys_tmp3773;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h39)) begin
										r_sub08_result_datain <= w_sys_tmp3855;

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3a)) begin
										r_sub08_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3a)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3b)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp2844[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_T_datain <= w_sys_tmp2847;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp2836[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_V_datain <= w_sys_tmp2839;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp2828[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_U_datain <= w_sys_tmp2831;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h6f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub12_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp3811[14:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp3820[14:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp3894[14:0] );

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h3d)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp3899[14:0] );

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp6806[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub12_result_datain <= w_sys_tmp3813;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h3d)) begin
										r_sub12_result_datain <= w_sys_tmp3903;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h3d)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp897[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_T_datain <= w_sys_tmp900;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp889[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_V_datain <= w_sys_tmp892;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp881[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_U_datain <= w_sys_tmp884;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub03_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3697[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp3694[14:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp5259[14:0] );

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp5248[14:0] );

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp5971[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub03_result_datain <= w_sys_tmp3721;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub03_result_datain <= w_sys_tmp5252;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hd6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp682[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_T_datain <= w_sys_tmp685;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp674[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_V_datain <= w_sys_tmp677;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp666[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_U_datain <= w_sys_tmp669;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3697[14:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3703[14:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3691[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp3694[14:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp4801[14:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp4812[14:0] );

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp5875[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub02_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub02_result_datain <= w_sys_tmp3693;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub02_result_datain <= w_sys_tmp4805;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hd0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp2625[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_T_datain <= w_sys_tmp2628;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp2617[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_V_datain <= w_sys_tmp2620;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp2609[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_U_datain <= w_sys_tmp2612;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h64: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub11_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3777[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp3774[14:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5289[14:0] );

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5279[14:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5273[14:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h59)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp5299[14:0] );

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp6707[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub11_result_datain <= w_sys_tmp3801;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub11_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub11_result_datain <= w_sys_tmp5252;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h57) || (r_sys_run_step==7'h58)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h59)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3274[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_T_datain <= w_sys_tmp3277;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp3266[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_V_datain <= w_sys_tmp3269;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp3258[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_U_datain <= w_sys_tmp3261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub14_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp3823[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp3814[14:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp3817[14:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp3842[14:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4846[14:0] );

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4852[14:0] );

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp4842[14:0] );

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp6979[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sub14_result_datain <= w_sys_tmp3813;

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub14_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub14_result_datain <= w_sys_tmp4856;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp467[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_T_datain <= w_sys_tmp470;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp459[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_V_datain <= w_sys_tmp462;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp451[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_U_datain <= w_sys_tmp454;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub01_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3697[14:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3703[14:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3691[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3694[14:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp4354[14:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp4365[14:0] );

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp5779[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub01_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub01_result_datain <= w_sys_tmp3699;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub01_result_datain <= w_sys_tmp4358;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3059[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_T_datain <= w_sys_tmp3062;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp3051[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_V_datain <= w_sys_tmp3054;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp3043[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_U_datain <= w_sys_tmp3046;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h75: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub13_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp3811[14:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp3823[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp3814[14:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp3817[14:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4399[14:0] );

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4395[14:0] );

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp4405[14:0] );

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp6883[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub13_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub13_result_datain <= w_sys_tmp3819;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub13_result_datain <= w_sys_tmp4409;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp252[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_T_datain <= w_sys_tmp255;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp244[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_V_datain <= w_sys_tmp247;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp236[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_U_datain <= w_sys_tmp239;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub00_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3700[14:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3691[14:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3851[14:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3866[14:0] );

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp5702[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_datain <= w_sys_tmp3693;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32)) begin
										r_sub00_result_datain <= w_sys_tmp3855;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h32)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hc4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp1761[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_T_datain <= w_sys_tmp1764;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1753[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_V_datain <= w_sys_tmp1756;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1745[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_U_datain <= w_sys_tmp1748;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub07_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3737[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3734[14:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp5259[14:0] );

									end
									else
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h55)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp5279[14:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp5253[14:0] );

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp5269[14:0] );

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp6339[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub07_result_datain <= w_sys_tmp3761;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub07_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub07_result_datain <= w_sys_tmp5263;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h53) || (r_sys_run_step==7'h54)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h55)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hf3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp1546[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_T_datain <= w_sys_tmp1549;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1538[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_V_datain <= w_sys_tmp1541;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1530[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_U_datain <= w_sys_tmp1533;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub06_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3731[14:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3743[14:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3737[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3734[14:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4806[14:0] );

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4822[14:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4812[14:0] );

									end
									else
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h55)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp4832[14:0] );

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp6243[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub06_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_result_datain <= w_sys_tmp3733;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub06_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub06_result_datain <= w_sys_tmp4816;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h53) || (r_sys_run_step==7'h54)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h55)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3489[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_T_datain <= w_sys_tmp3492;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp3481[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_V_datain <= w_sys_tmp3484;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp3473[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_U_datain <= w_sys_tmp3476;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h81: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub15_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3814[14:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp3817[14:0] );

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5293[14:0] );

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5289[14:0] );

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp5299[14:0] );

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp7075[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub15_result_datain <= w_sys_tmp3841;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub15_result_datain <= w_sys_tmp5303;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h5b)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h42) || (r_sys_run_step==7'h4f)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp1331[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_T_datain <= w_sys_tmp1334;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1323[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_V_datain <= w_sys_tmp1326;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1315[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_U_datain <= w_sys_tmp1318;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h3b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3731[14:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3743[14:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3737[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3734[14:0] );

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4359[14:0] );

									end
									else
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h55)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4385[14:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4365[14:0] );

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp4375[14:0] );

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp6147[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub05_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub05_result_datain <= w_sys_tmp3739;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h54)) begin
										r_sub05_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h53)) begin
										r_sub05_result_datain <= w_sys_tmp4369;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h3a) || (r_sys_run_step==7'h46) || (r_sys_run_step==7'h47) || (r_sys_run_step==7'h53) || (r_sys_run_step==7'h54)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h48) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h55)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1116[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_T_datain <= w_sys_tmp1119;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1108[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_V_datain <= w_sys_tmp1111;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1100[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_U_datain <= w_sys_tmp1103;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h35: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub04_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3740[14:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3731[14:0] );

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3861[14:0] );

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3871[14:0] );

									end
									else
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h37)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3885[14:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h30)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp3856[14:0] );

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp6070[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_datain <= w_sys_tmp3733;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h35)) begin
										r_sub04_result_datain <= w_sys_tmp3865;

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub04_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h36)) begin
										r_sub04_result_datain <= w_sys_tmp3903;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h36)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h37)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp2410[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_T_datain <= w_sys_tmp2413;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp2402[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_V_datain <= w_sys_tmp2405;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp2394[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_U_datain <= w_sys_tmp2397;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h5e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub10_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3783[14:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3777[14:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3771[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp3774[14:0] );

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h59)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4852[14:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4842[14:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4e)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4826[14:0] );

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4832[14:0] );

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp6611[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sub10_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub10_result_datain <= w_sys_tmp3773;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h58)) begin
										r_sub10_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h57)) begin
										r_sub10_result_datain <= w_sys_tmp4805;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'h87: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h4b) || (r_sys_run_step==7'h57) || (r_sys_run_step==7'h58)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h4c) || (r_sys_run_step==7'h4e) || (r_sys_run_step==7'h59)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						9'h12f: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp0_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp0_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp0_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sys_tmp0_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						9'h8f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						9'h95: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp1_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						9'h9b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp1_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						9'ha7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h38)) begin
										r_sys_tmp1_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sys_tmp1_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h12) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19)) begin
										r_sys_tmp2_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp2_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h50)) begin
										r_sys_tmp2_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						9'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sys_tmp2_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17)) begin
										r_sys_tmp3_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						9'ha1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp3_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						9'had: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sys_tmp3_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						9'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'hd)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==7'hf) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						9'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h44) || (r_sys_run_step==7'h51)) begin
										r_sys_tmp4_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
