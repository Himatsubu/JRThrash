/*
TimeStamp:	2016/12/20		15:43
*/


module NeuralNet(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_threadTop_req,	
	output                o_threadTop_busy	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg         [31:0] r_ip_DivFloat_dividend_0;
	reg         [31:0] r_ip_DivFloat_divisor_0;
	wire        [31:0] w_ip_DivFloat_quotient_0;
	reg         [31:0] r_ip_CompareFloatLT_portA_0;
	reg         [31:0] r_ip_CompareFloatLT_portB_0;
	wire               w_ip_CompareFloatLT_result_0;
	wire        [31:0] w_ip_rand_result_0;
	wire        [31:0] w_ip_rand_result_1;
	wire        [31:0] w_ip_rand_result_2;
	wire        [31:0] w_ip_rand_result_3;
	wire        [31:0] w_ip_rand_result_4;
	wire        [31:0] w_ip_rand_result_5;
	wire        [31:0] w_ip_rand_result_6;
	wire        [31:0] w_ip_rand_result_7;
	wire        [31:0] w_ip_rand_result_8;
	wire        [31:0] w_ip_rand_result_9;
	reg         [31:0] r_ip_exp_i_0;
	wire        [31:0] w_ip_exp_result_0;
	reg         [31:0] r_ip_exp_i_1;
	wire        [31:0] w_ip_exp_result_1;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_threadTop_caller;
	reg                r_sys_threadTop_req;
	reg         [ 6:0] r_sys_threadTop_phase;
	reg         [ 1:0] r_sys_threadTop_stage;
	reg         [ 6:0] r_sys_threadTop_step;
	reg                r_sys_threadTop_busy;
	wire        [ 1:0] w_sys_threadTop_stage_p1;
	wire        [ 6:0] w_sys_threadTop_step_p1;
	reg  signed [31:0] r_fld_N_INPUT_0;
	reg  signed [31:0] r_fld_N_HIDDEN_1;
	reg  signed [31:0] r_fld_N_OUTPUT_2;
	wire signed [ 3:0] w_fld_w1_3_addr_0;
	wire        [31:0] w_fld_w1_3_datain_0;
	wire        [31:0] w_fld_w1_3_dataout_0;
	wire               w_fld_w1_3_r_w_0;
	wire               w_fld_w1_3_ce_0;
	reg  signed [ 3:0] r_fld_w1_3_addr_1;
	reg         [31:0] r_fld_w1_3_datain_1;
	wire        [31:0] w_fld_w1_3_dataout_1;
	reg                r_fld_w1_3_r_w_1;
	wire               w_fld_w1_3_ce_1;
	wire signed [ 2:0] w_fld_w2_4_addr_0;
	wire        [31:0] w_fld_w2_4_datain_0;
	wire        [31:0] w_fld_w2_4_dataout_0;
	wire               w_fld_w2_4_r_w_0;
	wire               w_fld_w2_4_ce_0;
	reg  signed [ 2:0] r_fld_w2_4_addr_1;
	reg         [31:0] r_fld_w2_4_datain_1;
	wire        [31:0] w_fld_w2_4_dataout_1;
	reg                r_fld_w2_4_r_w_1;
	wire               w_fld_w2_4_ce_1;
	wire signed        w_fld_input_5_addr_0;
	wire        [31:0] w_fld_input_5_datain_0;
	wire        [31:0] w_fld_input_5_dataout_0;
	wire               w_fld_input_5_r_w_0;
	wire               w_fld_input_5_ce_0;
	reg  signed        r_fld_input_5_addr_1;
	reg         [31:0] r_fld_input_5_datain_1;
	wire        [31:0] w_fld_input_5_dataout_1;
	reg                r_fld_input_5_r_w_1;
	wire               w_fld_input_5_ce_1;
	wire signed [ 2:0] w_fld_hidden_6_addr_0;
	wire        [31:0] w_fld_hidden_6_datain_0;
	wire        [31:0] w_fld_hidden_6_dataout_0;
	wire               w_fld_hidden_6_r_w_0;
	wire               w_fld_hidden_6_ce_0;
	reg  signed [ 2:0] r_fld_hidden_6_addr_1;
	reg         [31:0] r_fld_hidden_6_datain_1;
	wire        [31:0] w_fld_hidden_6_dataout_1;
	reg                r_fld_hidden_6_r_w_1;
	wire               w_fld_hidden_6_ce_1;
	wire signed        w_fld_output_7_addr_0;
	wire        [31:0] w_fld_output_7_datain_0;
	wire        [31:0] w_fld_output_7_dataout_0;
	wire               w_fld_output_7_r_w_0;
	wire               w_fld_output_7_ce_0;
	reg  signed        r_fld_output_7_addr_1;
	reg         [31:0] r_fld_output_7_datain_1;
	wire        [31:0] w_fld_output_7_dataout_1;
	reg                r_fld_output_7_r_w_1;
	wire               w_fld_output_7_ce_1;
	wire signed [ 2:0] w_fld_in_8_addr_0;
	wire        [31:0] w_fld_in_8_datain_0;
	wire        [31:0] w_fld_in_8_dataout_0;
	wire               w_fld_in_8_r_w_0;
	wire               w_fld_in_8_ce_0;
	reg  signed [ 2:0] r_fld_in_8_addr_1;
	reg         [31:0] r_fld_in_8_datain_1;
	wire        [31:0] w_fld_in_8_dataout_1;
	reg                r_fld_in_8_r_w_1;
	wire               w_fld_in_8_ce_1;
	wire signed [ 1:0] w_fld_res_9_addr_0;
	wire        [31:0] w_fld_res_9_datain_0;
	wire        [31:0] w_fld_res_9_dataout_0;
	wire               w_fld_res_9_r_w_0;
	wire               w_fld_res_9_ce_0;
	reg  signed [ 1:0] r_fld_res_9_addr_1;
	reg         [31:0] r_fld_res_9_datain_1;
	wire        [31:0] w_fld_res_9_dataout_1;
	reg                r_fld_res_9_r_w_1;
	wire               w_fld_res_9_ce_1;
	reg         [31:0] r_threadTop_err_10;
	reg         [31:0] r_threadTop_alpha_11;
	reg         [31:0] r_threadTop_sum_12;
	reg         [31:0] r_threadTop_delta_13;
	reg  signed [31:0] r_threadTop_i_14;
	reg  signed [31:0] r_threadTop_j_15;
	reg  signed [31:0] r_threadTop_i_16;
	reg  signed [31:0] r_threadTop_j_17;
	reg  signed [31:0] r_threadTop_i_18;
	reg  signed [31:0] r_threadTop_j_19;
	reg  signed [31:0] r_threadTop_k_20;
	reg  signed [31:0] r_threadTop_j_21;
	reg  signed [31:0] r_threadTop_k_22;
	reg  signed [31:0] r_threadTop_j_23;
	reg  signed [31:0] r_threadTop_k_24;
	reg  signed [31:0] r_threadTop_j_25;
	reg  signed [31:0] r_threadTop_l_26;
	reg  signed [31:0] r_threadTop_k_27;
	reg  signed [31:0] r_threadTop_j_28;
	reg  signed [31:0] r_threadTop_k_29;
	reg  signed [31:0] r_threadTop_copy0_j_31;
	reg  signed [31:0] r_threadTop_copy0_j_32;
	reg  signed [31:0] r_threadTop_copy0_j_33;
	reg  signed [31:0] r_threadTop_copy0_j_34;
	reg  signed [31:0] r_threadTop_copy1_j_35;
	reg  signed [31:0] r_threadTop_copy0_j_36;
	reg  signed [31:0] r_threadTop_copy1_j_37;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	wire        [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire signed [31:0] w_sys_tmp7;
	wire signed [31:0] w_sys_tmp10;
	wire signed [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp22;
	wire               w_sys_tmp34;
	wire signed [31:0] w_sys_tmp35;
	wire               w_sys_tmp36;
	wire signed [31:0] w_sys_tmp39;
	wire signed [31:0] w_sys_tmp40;
	wire signed [31:0] w_sys_tmp41;
	wire        [31:0] w_sys_tmp42;
	wire        [31:0] w_sys_tmp43;
	wire        [31:0] w_sys_tmp45;
	wire        [31:0] w_sys_tmp46;
	wire        [31:0] w_sys_tmp47;
	wire        [31:0] w_sys_tmp48;
	wire signed [31:0] w_sys_tmp49;
	wire               w_sys_tmp94;
	wire signed [31:0] w_sys_tmp95;
	wire               w_sys_tmp96;
	wire signed [31:0] w_sys_tmp99;
	wire        [31:0] w_sys_tmp100;
	wire        [31:0] w_sys_tmp101;
	wire        [31:0] w_sys_tmp103;
	wire        [31:0] w_sys_tmp104;
	wire        [31:0] w_sys_tmp105;
	wire        [31:0] w_sys_tmp106;
	wire signed [31:0] w_sys_tmp107;
	wire        [31:0] w_sys_tmp144;
	wire               w_sys_tmp145;
	wire signed [31:0] w_sys_tmp146;
	wire               w_sys_tmp148;
	wire        [31:0] w_sys_tmp151;
	wire signed [31:0] w_sys_tmp152;
	wire signed [31:0] w_sys_tmp153;
	wire signed [31:0] w_sys_tmp154;
	wire signed [31:0] w_sys_tmp155;
	wire signed [31:0] w_sys_tmp156;
	wire               w_sys_tmp185;
	wire        [31:0] w_sys_tmp188;
	wire               w_sys_tmp189;
	wire        [31:0] w_sys_tmp192;
	wire        [31:0] w_sys_tmp193;
	wire        [31:0] w_sys_tmp194;
	wire signed [31:0] w_sys_tmp195;
	wire signed [31:0] w_sys_tmp196;
	wire signed [31:0] w_sys_tmp197;
	wire        [31:0] w_sys_tmp198;
	wire signed [31:0] w_sys_tmp199;
	wire signed [31:0] w_sys_tmp200;
	wire        [31:0] w_sys_tmp203;
	wire        [31:0] w_sys_tmp242;
	wire        [31:0] w_sys_tmp243;
	wire        [31:0] w_sys_tmp244;
	wire        [31:0] w_sys_tmp246;
	wire        [31:0] w_sys_tmp247;
	wire        [31:0] w_sys_tmp248;
	wire signed [31:0] w_sys_tmp249;
	wire               w_sys_tmp250;
	wire        [31:0] w_sys_tmp253;
	wire               w_sys_tmp254;
	wire        [31:0] w_sys_tmp257;
	wire        [31:0] w_sys_tmp258;
	wire        [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp260;
	wire        [31:0] w_sys_tmp261;
	wire signed [31:0] w_sys_tmp262;
	wire signed [31:0] w_sys_tmp263;
	wire        [31:0] w_sys_tmp266;
	wire        [31:0] w_sys_tmp297;
	wire        [31:0] w_sys_tmp298;
	wire        [31:0] w_sys_tmp299;
	wire        [31:0] w_sys_tmp301;
	wire        [31:0] w_sys_tmp302;
	wire        [31:0] w_sys_tmp303;
	wire signed [31:0] w_sys_tmp304;
	wire               w_sys_tmp305;
	wire signed [31:0] w_sys_tmp306;
	wire               w_sys_tmp307;
	wire        [31:0] w_sys_tmp309;
	wire        [31:0] w_sys_tmp310;
	wire        [31:0] w_sys_tmp314;
	wire        [31:0] w_sys_tmp315;
	wire        [31:0] w_sys_tmp316;
	wire signed [31:0] w_sys_tmp317;
	wire        [31:0] w_sys_tmp318;
	wire        [31:0] w_sys_tmp319;
	wire signed [31:0] w_sys_tmp322;
	wire signed [31:0] w_sys_tmp324;
	wire        [31:0] w_sys_tmp325;
	wire signed [31:0] w_sys_tmp326;
	wire signed [31:0] w_sys_tmp327;
	wire signed [31:0] w_sys_tmp328;
	wire        [31:0] w_sys_tmp343;
	wire               w_sys_tmp402;
	wire signed [31:0] w_sys_tmp403;
	wire        [31:0] w_sys_tmp404;
	wire               w_sys_tmp405;
	wire        [31:0] w_sys_tmp407;
	wire        [31:0] w_sys_tmp408;
	wire signed [31:0] w_sys_tmp411;
	wire        [31:0] w_sys_tmp413;
	wire signed [31:0] w_sys_tmp414;
	wire        [31:0] w_sys_tmp415;
	wire        [31:0] w_sys_tmp416;
	wire signed [31:0] w_sys_tmp418;
	wire               w_sys_tmp419;
	wire        [31:0] w_sys_tmp421;
	wire        [31:0] w_sys_tmp424;
	wire        [31:0] w_sys_tmp425;
	wire        [31:0] w_sys_tmp426;
	wire signed [31:0] w_sys_tmp429;
	wire signed [31:0] w_sys_tmp430;
	wire signed [31:0] w_sys_tmp431;
	wire signed [31:0] w_sys_tmp433;
	wire signed [31:0] w_sys_tmp434;
	wire        [31:0] w_sys_tmp436;
	wire signed [31:0] w_sys_tmp437;
	wire signed [31:0] w_sys_tmp438;
	wire signed [31:0] w_sys_tmp439;
	wire        [31:0] w_sys_tmp452;
	wire        [31:0] w_sys_tmp513;
	wire               w_sys_tmp514;
	wire        [31:0] w_sys_tmp516;
	wire        [31:0] w_sys_tmp517;
	wire        [31:0] w_sys_tmp518;
	wire signed [31:0] w_sys_tmp519;
	wire        [31:0] w_sys_tmp520;
	wire signed [31:0] w_sys_tmp525;
	wire        [31:0] w_sys_tmp526;
	wire        [31:0] w_sys_tmp527;
	wire signed [31:0] w_sys_tmp528;
	wire               w_sys_tmp529;
	wire        [31:0] w_sys_tmp530;
	wire signed [31:0] w_sys_tmp531;
	wire signed [31:0] w_sys_tmp532;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_threadTop_busy = r_sys_threadTop_busy;
	assign w_sys_threadTop_stage_p1 = (r_sys_threadTop_stage + 2'h1);
	assign w_sys_threadTop_step_p1 = (r_sys_threadTop_step + 7'h1);
	assign w_fld_w1_3_addr_0 = 4'sh0;
	assign w_fld_w1_3_datain_0 = 32'h0;
	assign w_fld_w1_3_r_w_0 = 1'h0;
	assign w_fld_w1_3_ce_0 = w_sys_ce;
	assign w_fld_w1_3_ce_1 = w_sys_ce;
	assign w_fld_w2_4_addr_0 = 3'sh0;
	assign w_fld_w2_4_datain_0 = 32'h0;
	assign w_fld_w2_4_r_w_0 = 1'h0;
	assign w_fld_w2_4_ce_0 = w_sys_ce;
	assign w_fld_w2_4_ce_1 = w_sys_ce;
	assign w_fld_input_5_addr_0 = 1'sh0;
	assign w_fld_input_5_datain_0 = 32'h0;
	assign w_fld_input_5_r_w_0 = 1'h0;
	assign w_fld_input_5_ce_0 = w_sys_ce;
	assign w_fld_input_5_ce_1 = w_sys_ce;
	assign w_fld_hidden_6_addr_0 = 3'sh0;
	assign w_fld_hidden_6_datain_0 = 32'h0;
	assign w_fld_hidden_6_r_w_0 = 1'h0;
	assign w_fld_hidden_6_ce_0 = w_sys_ce;
	assign w_fld_hidden_6_ce_1 = w_sys_ce;
	assign w_fld_output_7_addr_0 = 1'sh0;
	assign w_fld_output_7_datain_0 = 32'h0;
	assign w_fld_output_7_r_w_0 = 1'h0;
	assign w_fld_output_7_ce_0 = w_sys_ce;
	assign w_fld_output_7_ce_1 = w_sys_ce;
	assign w_fld_in_8_addr_0 = 3'sh0;
	assign w_fld_in_8_datain_0 = 32'h0;
	assign w_fld_in_8_r_w_0 = 1'h0;
	assign w_fld_in_8_ce_0 = w_sys_ce;
	assign w_fld_in_8_ce_1 = w_sys_ce;
	assign w_fld_res_9_addr_0 = 2'sh0;
	assign w_fld_res_9_datain_0 = 32'h0;
	assign w_fld_res_9_r_w_0 = 1'h0;
	assign w_fld_res_9_ce_0 = w_sys_ce;
	assign w_fld_res_9_ce_1 = w_sys_ce;
	assign w_sys_tmp1 = 32'h0;
	assign w_sys_tmp3 = 32'h3f800000;
	assign w_sys_tmp7 = 32'sh00000002;
	assign w_sys_tmp10 = 32'sh00000003;
	assign w_sys_tmp13 = 32'sh00000004;
	assign w_sys_tmp16 = 32'sh00000005;
	assign w_sys_tmp19 = 32'sh00000006;
	assign w_sys_tmp22 = 32'sh00000007;
	assign w_sys_tmp34 = (r_threadTop_i_14 < r_fld_N_INPUT_0);
	assign w_sys_tmp35 = (r_threadTop_i_14 + w_sys_intOne);
	assign w_sys_tmp36 = (r_threadTop_j_15 < r_fld_N_HIDDEN_1);
	assign w_sys_tmp39 = (w_sys_tmp40 + r_threadTop_j_15);
	assign w_sys_tmp40 = (w_sys_tmp41 * r_threadTop_i_14);
	assign w_sys_tmp41 = 32'sh00000005;
	assign w_sys_tmp42 = w_ip_MultFloat_product_0;
	assign w_sys_tmp43 = w_ip_AddFloat_result_0;
	assign w_sys_tmp45 = w_ip_rand_result_0;
	assign w_sys_tmp46 = 32'h40000000;
	assign w_sys_tmp47 = 32'h3f800000;
	assign w_sys_tmp48 = 32'h3dcccccd;
	assign w_sys_tmp49 = (r_threadTop_j_15 + w_sys_intOne);
	assign w_sys_tmp94 = (r_threadTop_i_16 < r_fld_N_HIDDEN_1);
	assign w_sys_tmp95 = (r_threadTop_i_16 + w_sys_intOne);
	assign w_sys_tmp96 = (r_threadTop_j_17 < r_fld_N_OUTPUT_2);
	assign w_sys_tmp99 = (r_threadTop_i_16 + r_threadTop_j_17);
	assign w_sys_tmp100 = w_ip_MultFloat_product_0;
	assign w_sys_tmp101 = w_ip_AddFloat_result_0;
	assign w_sys_tmp103 = w_ip_rand_result_5;
	assign w_sys_tmp104 = 32'h40000000;
	assign w_sys_tmp105 = 32'h3f800000;
	assign w_sys_tmp106 = 32'h3dcccccd;
	assign w_sys_tmp107 = (r_threadTop_j_17 + w_sys_intOne);
	assign w_sys_tmp144 = 32'h3dcccccd;
	assign w_sys_tmp145 = (r_threadTop_i_18 < w_sys_tmp146);
	assign w_sys_tmp146 = 32'sh00000004;
	assign w_sys_tmp148 = (r_threadTop_j_19 < r_fld_N_INPUT_0);
	assign w_sys_tmp151 = w_fld_in_8_dataout_1;
	assign w_sys_tmp152 = (w_sys_tmp153 + r_threadTop_copy0_j_31);
	assign w_sys_tmp153 = (w_sys_tmp154 * r_threadTop_i_18);
	assign w_sys_tmp154 = 32'sh00000002;
	assign w_sys_tmp155 = (r_threadTop_copy0_j_31 + w_sys_intOne);
	assign w_sys_tmp156 = (r_threadTop_j_19 + w_sys_intOne);
	assign w_sys_tmp185 = (r_threadTop_k_20 < r_fld_N_HIDDEN_1);
	assign w_sys_tmp188 = 32'h0;
	assign w_sys_tmp189 = (r_threadTop_j_21 < r_fld_N_INPUT_0);
	assign w_sys_tmp192 = w_ip_AddFloat_result_0;
	assign w_sys_tmp193 = w_ip_MultFloat_product_0;
	assign w_sys_tmp194 = w_fld_w1_3_dataout_1;
	assign w_sys_tmp195 = (w_sys_tmp196 + r_threadTop_k_20);
	assign w_sys_tmp196 = (w_sys_tmp197 * r_threadTop_j_21);
	assign w_sys_tmp197 = 32'sh00000005;
	assign w_sys_tmp198 = w_fld_input_5_dataout_1;
	assign w_sys_tmp199 = (r_threadTop_copy0_j_32 + w_sys_intOne);
	assign w_sys_tmp200 = (r_threadTop_j_21 + w_sys_intOne);
	assign w_sys_tmp203 = w_fld_hidden_6_dataout_1;
	assign w_sys_tmp242 = w_ip_DivFloat_quotient_0;
	assign w_sys_tmp243 = 32'h3f800000;
	assign w_sys_tmp244 = w_ip_AddFloat_result_0;
	assign w_sys_tmp246 = w_ip_exp_result_0;
	assign w_sys_tmp247 = ( -w_sys_tmp248 );
	assign w_sys_tmp248 = w_fld_hidden_6_dataout_1;
	assign w_sys_tmp249 = (r_threadTop_k_20 + w_sys_intOne);
	assign w_sys_tmp250 = (r_threadTop_k_22 < r_fld_N_OUTPUT_2);
	assign w_sys_tmp253 = 32'h0;
	assign w_sys_tmp254 = (r_threadTop_j_23 < r_fld_N_HIDDEN_1);
	assign w_sys_tmp257 = w_ip_AddFloat_result_0;
	assign w_sys_tmp258 = w_ip_MultFloat_product_0;
	assign w_sys_tmp259 = w_fld_w2_4_dataout_1;
	assign w_sys_tmp260 = (r_threadTop_j_23 + r_threadTop_k_22);
	assign w_sys_tmp261 = w_fld_hidden_6_dataout_1;
	assign w_sys_tmp262 = (r_threadTop_copy0_j_33 + w_sys_intOne);
	assign w_sys_tmp263 = (r_threadTop_j_23 + w_sys_intOne);
	assign w_sys_tmp266 = w_fld_output_7_dataout_1;
	assign w_sys_tmp297 = w_ip_DivFloat_quotient_0;
	assign w_sys_tmp298 = 32'h3f800000;
	assign w_sys_tmp299 = w_ip_AddFloat_result_0;
	assign w_sys_tmp301 = w_ip_exp_result_1;
	assign w_sys_tmp302 = ( -w_sys_tmp303 );
	assign w_sys_tmp303 = w_fld_output_7_dataout_1;
	assign w_sys_tmp304 = (r_threadTop_k_22 + w_sys_intOne);
	assign w_sys_tmp305 = (r_threadTop_k_24 < r_fld_N_OUTPUT_2);
	assign w_sys_tmp306 = (r_threadTop_k_24 + w_sys_intOne);
	assign w_sys_tmp307 = (r_threadTop_j_25 < r_fld_N_HIDDEN_1);
	assign w_sys_tmp309 = w_ip_MultFloat_product_0;
	assign w_sys_tmp310 = ( -r_threadTop_alpha_11 );
	assign w_sys_tmp314 = ( -w_sys_tmp315 );
	assign w_sys_tmp315 = w_ip_AddFloat_result_0;
	assign w_sys_tmp316 = w_fld_res_9_dataout_1;
	assign w_sys_tmp317 = (r_threadTop_i_18 + r_threadTop_k_24);
	assign w_sys_tmp318 = w_fld_output_7_dataout_1;
	assign w_sys_tmp319 = 32'h3f800000;
	assign w_sys_tmp322 = (r_threadTop_copy1_j_35 + r_threadTop_k_24);
	assign w_sys_tmp324 = (r_threadTop_copy0_j_34 + r_threadTop_k_24);
	assign w_sys_tmp325 = w_sys_tmp309;
	assign w_sys_tmp326 = (r_threadTop_copy0_j_34 + w_sys_intOne);
	assign w_sys_tmp327 = (r_threadTop_copy1_j_35 + w_sys_intOne);
	assign w_sys_tmp328 = (r_threadTop_j_25 + w_sys_intOne);
	assign w_sys_tmp343 = w_fld_w2_4_dataout_1;
	assign w_sys_tmp402 = (r_threadTop_l_26 < r_fld_N_HIDDEN_1);
	assign w_sys_tmp403 = (r_threadTop_l_26 + w_sys_intOne);
	assign w_sys_tmp404 = 32'h0;
	assign w_sys_tmp405 = (r_threadTop_k_27 < r_fld_N_OUTPUT_2);
	assign w_sys_tmp407 = w_ip_AddFloat_result_0;
	assign w_sys_tmp408 = w_ip_MultFloat_product_0;
	assign w_sys_tmp411 = (r_threadTop_l_26 + r_threadTop_k_27);
	assign w_sys_tmp413 = w_fld_res_9_dataout_1;
	assign w_sys_tmp414 = (r_threadTop_i_18 + r_threadTop_k_27);
	assign w_sys_tmp415 = w_fld_output_7_dataout_1;
	assign w_sys_tmp416 = 32'h3f800000;
	assign w_sys_tmp418 = (r_threadTop_k_27 + w_sys_intOne);
	assign w_sys_tmp419 = (r_threadTop_j_28 < r_fld_N_INPUT_0);
	assign w_sys_tmp421 = w_ip_MultFloat_product_0;
	assign w_sys_tmp424 = w_fld_hidden_6_dataout_1;
	assign w_sys_tmp425 = w_ip_AddFloat_result_0;
	assign w_sys_tmp426 = 32'h3f800000;
	assign w_sys_tmp429 = (w_sys_tmp430 + r_threadTop_l_26);
	assign w_sys_tmp430 = (w_sys_tmp431 * r_threadTop_copy1_j_37);
	assign w_sys_tmp431 = 32'sh00000005;
	assign w_sys_tmp433 = (w_sys_tmp434 + r_threadTop_l_26);
	assign w_sys_tmp434 = (w_sys_tmp431 * r_threadTop_copy0_j_36);
	assign w_sys_tmp436 = w_sys_tmp421;
	assign w_sys_tmp437 = (r_threadTop_copy0_j_36 + w_sys_intOne);
	assign w_sys_tmp438 = (r_threadTop_copy1_j_37 + w_sys_intOne);
	assign w_sys_tmp439 = (r_threadTop_j_28 + w_sys_intOne);
	assign w_sys_tmp452 = w_fld_w1_3_dataout_1;
	assign w_sys_tmp513 = 32'h0;
	assign w_sys_tmp514 = (r_threadTop_k_29 < r_fld_N_OUTPUT_2);
	assign w_sys_tmp516 = w_ip_AddFloat_result_0;
	assign w_sys_tmp517 = w_ip_MultFloat_product_0;
	assign w_sys_tmp518 = w_fld_res_9_dataout_1;
	assign w_sys_tmp519 = (r_threadTop_i_18 + r_threadTop_k_29);
	assign w_sys_tmp520 = w_fld_output_7_dataout_1;
	assign w_sys_tmp525 = (r_threadTop_k_29 + w_sys_intOne);
	assign w_sys_tmp526 = w_ip_MultFloat_product_0;
	assign w_sys_tmp527 = 32'h3f000000;
	assign w_sys_tmp528 = (r_threadTop_i_18 + w_sys_intOne);
	assign w_sys_tmp529 = w_ip_CompareFloatLT_result_0;
	assign w_sys_tmp530 = 32'h3a83126f;
	assign w_sys_tmp531 = 32'sh00000002;
	assign w_sys_tmp532 = 32'sh00000005;


	DualPortRAM #(.DWIDTH(32), .AWIDTH(4), .WORDS(10) )
		dpram_w1_3(
			.clk (clock),
			.ce_0 (w_fld_w1_3_ce_0),
			.addr_0 (w_fld_w1_3_addr_0),
			.datain_0 (w_fld_w1_3_datain_0),
			.dataout_0 (w_fld_w1_3_dataout_0),
			.r_w_0 (w_fld_w1_3_r_w_0),
			.ce_1 (w_fld_w1_3_ce_1),
			.addr_1 (r_fld_w1_3_addr_1),
			.datain_1 (r_fld_w1_3_datain_1),
			.dataout_1 (w_fld_w1_3_dataout_1),
			.r_w_1 (r_fld_w1_3_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(3), .WORDS(5) )
		dpram_w2_4(
			.clk (clock),
			.ce_0 (w_fld_w2_4_ce_0),
			.addr_0 (w_fld_w2_4_addr_0),
			.datain_0 (w_fld_w2_4_datain_0),
			.dataout_0 (w_fld_w2_4_dataout_0),
			.r_w_0 (w_fld_w2_4_r_w_0),
			.ce_1 (w_fld_w2_4_ce_1),
			.addr_1 (r_fld_w2_4_addr_1),
			.datain_1 (r_fld_w2_4_datain_1),
			.dataout_1 (w_fld_w2_4_dataout_1),
			.r_w_1 (r_fld_w2_4_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(1), .WORDS(2) )
		dpram_input_5(
			.clk (clock),
			.ce_0 (w_fld_input_5_ce_0),
			.addr_0 (w_fld_input_5_addr_0),
			.datain_0 (w_fld_input_5_datain_0),
			.dataout_0 (w_fld_input_5_dataout_0),
			.r_w_0 (w_fld_input_5_r_w_0),
			.ce_1 (w_fld_input_5_ce_1),
			.addr_1 (r_fld_input_5_addr_1),
			.datain_1 (r_fld_input_5_datain_1),
			.dataout_1 (w_fld_input_5_dataout_1),
			.r_w_1 (r_fld_input_5_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(3), .WORDS(5) )
		dpram_hidden_6(
			.clk (clock),
			.ce_0 (w_fld_hidden_6_ce_0),
			.addr_0 (w_fld_hidden_6_addr_0),
			.datain_0 (w_fld_hidden_6_datain_0),
			.dataout_0 (w_fld_hidden_6_dataout_0),
			.r_w_0 (w_fld_hidden_6_r_w_0),
			.ce_1 (w_fld_hidden_6_ce_1),
			.addr_1 (r_fld_hidden_6_addr_1),
			.datain_1 (r_fld_hidden_6_datain_1),
			.dataout_1 (w_fld_hidden_6_dataout_1),
			.r_w_1 (r_fld_hidden_6_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(1), .WORDS(1) )
		dpram_output_7(
			.clk (clock),
			.ce_0 (w_fld_output_7_ce_0),
			.addr_0 (w_fld_output_7_addr_0),
			.datain_0 (w_fld_output_7_datain_0),
			.dataout_0 (w_fld_output_7_dataout_0),
			.r_w_0 (w_fld_output_7_r_w_0),
			.ce_1 (w_fld_output_7_ce_1),
			.addr_1 (r_fld_output_7_addr_1),
			.datain_1 (r_fld_output_7_datain_1),
			.dataout_1 (w_fld_output_7_dataout_1),
			.r_w_1 (r_fld_output_7_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(3), .WORDS(8) )
		dpram_in_8(
			.clk (clock),
			.ce_0 (w_fld_in_8_ce_0),
			.addr_0 (w_fld_in_8_addr_0),
			.datain_0 (w_fld_in_8_datain_0),
			.dataout_0 (w_fld_in_8_dataout_0),
			.r_w_0 (w_fld_in_8_r_w_0),
			.ce_1 (w_fld_in_8_ce_1),
			.addr_1 (r_fld_in_8_addr_1),
			.datain_1 (r_fld_in_8_datain_1),
			.dataout_1 (w_fld_in_8_dataout_1),
			.r_w_1 (r_fld_in_8_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(2), .WORDS(4) )
		dpram_res_9(
			.clk (clock),
			.ce_0 (w_fld_res_9_ce_0),
			.addr_0 (w_fld_res_9_addr_0),
			.datain_0 (w_fld_res_9_datain_0),
			.dataout_0 (w_fld_res_9_dataout_0),
			.r_w_0 (w_fld_res_9_r_w_0),
			.ce_1 (w_fld_res_9_ce_1),
			.addr_1 (r_fld_res_9_addr_1),
			.datain_1 (r_fld_res_9_datain_1),
			.dataout_1 (w_fld_res_9_dataout_1),
			.r_w_1 (r_fld_res_9_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	DivFloat
		DivFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_DivFloat_dividend_0),
			.b (r_ip_DivFloat_divisor_0),
			.result (w_ip_DivFloat_quotient_0)
		);

	CompareFloatLT
		CompareFloatLT_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_CompareFloatLT_portA_0),
			.b (r_ip_CompareFloatLT_portB_0),
			.result (w_ip_CompareFloatLT_result_0)
		);

	rand
		rand_inst_0(
			.out (w_ip_rand_result_0)	// out 32bit
		);

	rand
		rand_inst_1(
			.out (w_ip_rand_result_1)	// out 32bit
		);

	rand
		rand_inst_2(
			.out (w_ip_rand_result_2)	// out 32bit
		);

	rand
		rand_inst_3(
			.out (w_ip_rand_result_3)	// out 32bit
		);

	rand
		rand_inst_4(
			.out (w_ip_rand_result_4)	// out 32bit
		);

	rand
		rand_inst_5(
			.out (w_ip_rand_result_5)	// out 32bit
		);

	rand
		rand_inst_6(
			.out (w_ip_rand_result_6)	// out 32bit
		);

	rand
		rand_inst_7(
			.out (w_ip_rand_result_7)	// out 32bit
		);

	rand
		rand_inst_8(
			.out (w_ip_rand_result_8)	// out 32bit
		);

	rand
		rand_inst_9(
			.out (w_ip_rand_result_9)	// out 32bit
		);

	exp
		exp_inst_0(
			.i (r_ip_exp_i_0),	// in 32bit
			.out (w_ip_exp_result_0)	// out 32bit
		);

	exp
		exp_inst_1(
			.i (r_ip_exp_i_1),	// in 32bit
			.out (w_ip_exp_result_1)	// out 32bit
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h5<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h9)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp42;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h5<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h9)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp100;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hf) || (r_sys_threadTop_step==7'h17) || (r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h27)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp203;

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp3_float;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp243;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_threadTop_step==7'hf) || (r_sys_threadTop_step==7'h17) || (r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h27)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp266;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp298;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_threadTop_step==7'h5) || (r_sys_threadTop_step==7'hb)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_threadTop_step==7'h23) || (r_sys_threadTop_step==7'h2b) || (r_sys_threadTop_step==7'h33) || (r_sys_threadTop_step==7'h3b)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp343;

									end
									else
									if((r_sys_threadTop_step==7'h4) || (r_sys_threadTop_step==7'h7) || (r_sys_threadTop_step==7'ha) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h10)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp319;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp316;

									end
									else
									if((r_sys_threadTop_step==7'he)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp413;

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp416;

									end
									else
									if((r_sys_threadTop_step==7'h16)) begin
										r_ip_AddFloat_portA_0 <= r_threadTop_sum_12;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3) || (r_sys_threadTop_step==7'h5) || (r_sys_threadTop_step==7'h7) || (r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hb)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp426;

									end
									else
									if((r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h27) || (r_sys_threadTop_step==7'h2f) || (r_sys_threadTop_step==7'h37)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp452;

									end
									else
									if((r_sys_threadTop_step==7'h17)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hd)) begin
										r_ip_AddFloat_portA_0 <= r_threadTop_err_10;

									end
									else
									if((r_sys_threadTop_step==7'h2) || (r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp518;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp47[31], w_sys_tmp47[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h9)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp47[31], w_sys_tmp47[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp47[31], w_sys_tmp47[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp47[31], w_sys_tmp47[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h5)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp47[31], w_sys_tmp47[30:0] };

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp105[31], w_sys_tmp105[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h9)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp105[31], w_sys_tmp105[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h6)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp105[31], w_sys_tmp105[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp105[31], w_sys_tmp105[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h5)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp105[31], w_sys_tmp105[30:0] };

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hf)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'h17)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp193;

									end
									else
									if((r_sys_threadTop_step==7'h27)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_threadTop_step==7'h1f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp246;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hf)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'h17)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_threadTop_step==7'h27)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_threadTop_step==7'h1f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp258;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp301;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hb)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp318[31], w_sys_tmp318[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'ha)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp318[31], w_sys_tmp318[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp318[31], w_sys_tmp318[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h1b)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp325;

									end
									else
									if((r_sys_threadTop_step==7'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp318[31], w_sys_tmp318[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp318[31], w_sys_tmp318[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h5)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp318[31], w_sys_tmp318[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp318[31], w_sys_tmp318[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp318[31], w_sys_tmp318[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp318[31], w_sys_tmp318[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h23) || (r_sys_threadTop_step==7'h2b) || (r_sys_threadTop_step==7'h33) || (r_sys_threadTop_step==7'h3b)) begin
										r_ip_AddFloat_portB_0 <= r_threadTop_delta_13;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp318[31], w_sys_tmp318[30:0] };

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h16)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp408;

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp415[31], w_sys_tmp415[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp415[31], w_sys_tmp415[30:0] };

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h17)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp436;

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp424[31], w_sys_tmp424[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp424[31], w_sys_tmp424[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h5)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp424[31], w_sys_tmp424[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h9)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp424[31], w_sys_tmp424[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h27) || (r_sys_threadTop_step==7'h2f) || (r_sys_threadTop_step==7'h37)) begin
										r_ip_AddFloat_portB_0 <= r_threadTop_delta_13;

									end
									else
									if((r_sys_threadTop_step==7'hb)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp424[31], w_sys_tmp424[30:0] };

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hd)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp517;

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp520[31], w_sys_tmp520[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp520[31], w_sys_tmp520[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'ha<=r_sys_threadTop_step && r_sys_threadTop_step<=7'he)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp43;

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp45;

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp103;

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp3_float;

									end
									else
									if((7'ha<=r_sys_threadTop_step && r_sys_threadTop_step<=7'he)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp101;

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp194;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp259;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7) || (r_sys_threadTop_step==7'ha) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h10) || (r_sys_threadTop_step==7'h13)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp314;

									end
									else
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'hf) || (r_sys_threadTop_step==7'h11) || (r_sys_threadTop_step==7'h12) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h17) || (r_sys_threadTop_step==7'h18) || (r_sys_threadTop_step==7'h1a) || (r_sys_threadTop_step==7'h1d)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp309;

									end
									else
									if((r_sys_threadTop_step==7'h16) || (r_sys_threadTop_step==7'h19) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h22)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp310;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'h11)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp408;

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2) || (r_sys_threadTop_step==7'h4) || (r_sys_threadTop_step==7'h6) || (r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hb)) begin
										r_ip_MultFloat_multiplicand_0 <= r_threadTop_alpha_11;

									end
									else
									if((7'hd<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h16) || (r_sys_threadTop_step==7'h18) || (r_sys_threadTop_step==7'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp421;

									end
									else
									if((r_sys_threadTop_step==7'h8) || (r_sys_threadTop_step==7'ha) || (r_sys_threadTop_step==7'hc)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp6_float;

									end
								end

							endcase
						end

						7'h66: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_ip_MultFloat_multiplicand_0 <= r_threadTop_err_10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'ha<=r_sys_threadTop_step && r_sys_threadTop_step<=7'he)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp48;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp46;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp104;

									end
									else
									if((7'ha<=r_sys_threadTop_step && r_sys_threadTop_step<=7'he)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp106;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp198;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp261;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'h1d)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_threadTop_step==7'ha) || (r_sys_threadTop_step==7'h10)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_threadTop_step==7'h7) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h13)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_threadTop_step==7'h17)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'hf) || (r_sys_threadTop_step==7'h12) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h18)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_threadTop_step==7'h11)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_threadTop_step==7'h16) || (r_sys_threadTop_step==7'h19) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h22)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp309;

									end
									else
									if((r_sys_threadTop_step==7'h14)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h11)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_threadTop_step==7'hc)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp407;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h13)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_threadTop_step==7'h2) || (r_sys_threadTop_step==7'h4) || (r_sys_threadTop_step==7'h6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp424;

									end
									else
									if((r_sys_threadTop_step==7'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_threadTop_step==7'h15)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_threadTop_step==7'hd)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_threadTop_step==7'h12) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h16) || (r_sys_threadTop_step==7'h18) || (r_sys_threadTop_step==7'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_threadTop_sum_12;

									end
									else
									if((r_sys_threadTop_step==7'h11)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_threadTop_step==7'h8) || (r_sys_threadTop_step==7'ha) || (r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'he) || (r_sys_threadTop_step==7'h10)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp425;

									end
									else
									if((r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hb)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp516;

									end
								end

							endcase
						end

						7'h66: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp527;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_DivFloat_dividend_0 <= w_sys_tmp243;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_DivFloat_dividend_0 <= w_sys_tmp298;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_DivFloat_divisor_0 <= w_sys_tmp244;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_DivFloat_divisor_0 <= w_sys_tmp299;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h68: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_ip_CompareFloatLT_portA_0 <= r_threadTop_err_10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h68: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_ip_CompareFloatLT_portB_0 <= w_sys_tmp530;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_exp_i_0 <= w_sys_tmp247;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_exp_i_1 <= w_sys_tmp302;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_threadTop_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h6c: begin
							r_sys_processing_methodID <= r_sys_threadTop_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h0: begin
							r_sys_threadTop_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7)) begin
										r_sys_threadTop_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp34) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp36) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h13)) begin
										r_sys_threadTop_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp94) ? 7'h14 : 7'h19);

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h15;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp96) ? 7'h18 : 7'h11);

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h13)) begin
										r_sys_threadTop_phase <= 7'h15;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h1b;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_boolFalse) ? 7'h1e : 7'h6c);

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h1f;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp145) ? 7'h23 : 7'h68);

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h24;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp148) ? 7'h27 : 7'h29);

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_threadTop_phase <= 7'h24;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h2a;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp185) ? 7'h2d : 7'h36);

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h2f;

									end
								end

							endcase
						end

						7'h2f: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h30;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp189) ? 7'h33 : 7'h34);

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_phase <= 7'h30;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_phase <= 7'h2a;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h37;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp250) ? 7'h3a : 7'h43);

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h3c;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h3d;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp254) ? 7'h40 : 7'h41);

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_phase <= 7'h3d;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_phase <= 7'h37;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h44;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp305) ? 7'h48 : 7'h4e);

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h44;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h49;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp307) ? 7'h4c : 7'h45);

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h40)) begin
										r_sys_threadTop_phase <= 7'h49;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h4f;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp402) ? 7'h52 : 7'h5f);

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h4f;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h54;

									end
								end

							endcase
						end

						7'h54: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h55;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp405) ? 7'h58 : 7'h5a);

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b)) begin
										r_sys_threadTop_phase <= 7'h55;

									end
								end

							endcase
						end

						7'h5a: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h5b;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp419) ? 7'h5e : 7'h50);

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3c)) begin
										r_sys_threadTop_phase <= 7'h5b;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h61;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h62;

									end
								end

							endcase
						end

						7'h62: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp514) ? 7'h65 : 7'h66);

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h12)) begin
										r_sys_threadTop_phase <= 7'h62;

									end
								end

							endcase
						end

						7'h66: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_sys_threadTop_phase <= 7'h1f;

									end
								end

							endcase
						end

						7'h68: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp529) ? 7'h6a : 7'h1b);

									end
								end

							endcase
						end

						7'h6a: begin
							r_sys_threadTop_phase <= 7'h6c;
						end

						7'h6c: begin
							r_sys_threadTop_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h13)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h13)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h40)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h54: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h5a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3c)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h62: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h12)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h66: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h68: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h13)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h12)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h14: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h12)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
									else
									if((r_sys_threadTop_step==7'h13)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h5)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h2b)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h25)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
									else
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h2b)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h25)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
									else
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h49: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3f)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
									else
									if((r_sys_threadTop_step==7'h40)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h52: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h54: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h55: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h1a)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h5a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h5b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3b)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
									else
									if((r_sys_threadTop_step==7'h3c)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h61: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h62: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h12)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h11)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h66: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
									else
									if((r_sys_threadTop_step==7'h5)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h68: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1) || (r_sys_threadTop_step==7'h2)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_threadTop_busy <= ((i_threadTop_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h0: begin
							r_sys_threadTop_busy <= w_sys_boolTrue;
						end

						7'h6c: begin
							r_sys_threadTop_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_N_INPUT_0 <= w_sys_tmp531;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_N_HIDDEN_1 <= w_sys_tmp532;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_N_OUTPUT_2 <= w_sys_intOne;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_w1_3_addr_1 <= 4'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'hf<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h13)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp39[3:0] );

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp195[3:0] );

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c) || (r_sys_threadTop_step==7'h34) || (r_sys_threadTop_step==7'h3c)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp429[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h25) || (r_sys_threadTop_step==7'h2d) || (r_sys_threadTop_step==7'h35)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp433[3:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'hf<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h13)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp42;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c) || (r_sys_threadTop_step==7'h34) || (r_sys_threadTop_step==7'h3c)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp425;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_w1_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'hf<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h13)) begin
										r_fld_w1_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_w1_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c) || (r_sys_threadTop_step==7'h34) || (r_sys_threadTop_step==7'h3c)) begin
										r_fld_w1_3_r_w_1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h25) || (r_sys_threadTop_step==7'h2d) || (r_sys_threadTop_step==7'h35)) begin
										r_fld_w1_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h6c: begin
							r_fld_w1_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_w2_4_addr_1 <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'hf<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h13)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp99[2:0] );

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp260[2:0] );

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h21) || (r_sys_threadTop_step==7'h29) || (r_sys_threadTop_step==7'h31) || (r_sys_threadTop_step==7'h39)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp324[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h20) || (r_sys_threadTop_step==7'h28) || (r_sys_threadTop_step==7'h30) || (r_sys_threadTop_step==7'h38) || (r_sys_threadTop_step==7'h40)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp322[2:0] );

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp411[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'hf<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h13)) begin
										r_fld_w2_4_datain_1 <= w_sys_tmp100;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h20) || (r_sys_threadTop_step==7'h28) || (r_sys_threadTop_step==7'h30) || (r_sys_threadTop_step==7'h38) || (r_sys_threadTop_step==7'h40)) begin
										r_fld_w2_4_datain_1 <= w_sys_tmp315;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_w2_4_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'hf<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h13)) begin
										r_fld_w2_4_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_w2_4_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h20) || (r_sys_threadTop_step==7'h28) || (r_sys_threadTop_step==7'h30) || (r_sys_threadTop_step==7'h38) || (r_sys_threadTop_step==7'h40)) begin
										r_fld_w2_4_r_w_1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h21) || (r_sys_threadTop_step==7'h29) || (r_sys_threadTop_step==7'h31) || (r_sys_threadTop_step==7'h39)) begin
										r_fld_w2_4_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w2_4_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h6c: begin
							r_fld_w2_4_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_input_5_addr_1 <= 1'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h27: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_fld_input_5_addr_1 <= $signed( r_threadTop_j_19[0:0] );

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_input_5_addr_1 <= $signed( r_threadTop_copy0_j_32[0:0] );

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_input_5_addr_1 <= $signed( r_threadTop_j_28[0:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h27: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_fld_input_5_datain_1 <= w_sys_tmp151;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_input_5_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h27: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_fld_input_5_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_input_5_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_input_5_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h6c: begin
							r_fld_input_5_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_hidden_6_addr_1 <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_k_20[2:0] );

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h25) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_k_20[2:0] );

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_i_18[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_k_20[2:0] );

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_copy0_j_33[2:0] );

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_j_25[2:0] );

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h9)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_l_26[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_datain_1 <= w_sys_tmp188;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_hidden_6_datain_1 <= w_sys_tmp192;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_hidden_6_datain_1 <= w_sys_tmp242;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h25)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h9)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h6c: begin
							r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_output_7_addr_1 <= 1'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h3a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_22[0:0] );

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h25) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_22[0:0] );

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h26)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_22[0:0] );

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'he)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_24[0:0] );

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1) || (r_sys_threadTop_step==7'h2)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_27[0:0] );

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_29[0:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h3a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_datain_1 <= w_sys_tmp253;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_output_7_datain_1 <= w_sys_tmp257;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_output_7_datain_1 <= w_sys_tmp297;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_output_7_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h3a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h25)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolTrue;

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'he)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1) || (r_sys_threadTop_step==7'h2)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h6c: begin
							r_fld_output_7_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_in_8_addr_1 <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp19[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h5)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp16[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp10[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_intZero[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_intOne[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp13[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp7[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp22[2:0] );

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp152[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1) || (r_sys_threadTop_step==7'h2) || (r_sys_threadTop_step==7'h5)) begin
										r_fld_in_8_datain_1 <= w_sys_tmp3;

									end
									else
									if((r_sys_threadTop_step==7'h3) || (r_sys_threadTop_step==7'h4) || (r_sys_threadTop_step==7'h6) || (r_sys_threadTop_step==7'h7)) begin
										r_fld_in_8_datain_1 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_in_8_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h7)) begin
										r_fld_in_8_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_in_8_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h6c: begin
							r_fld_in_8_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_res_9_addr_1 <= 2'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_tmp10[1:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_intZero[1:0] );

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_intOne[1:0] );

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_tmp7[1:0] );

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_tmp317[1:0] );

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_tmp414[1:0] );

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_tmp519[1:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1) || (r_sys_threadTop_step==7'h2)) begin
										r_fld_res_9_datain_1 <= w_sys_tmp3;

									end
									else
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h3)) begin
										r_fld_res_9_datain_1 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_res_9_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3)) begin
										r_fld_res_9_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_res_9_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_res_9_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1)) begin
										r_fld_res_9_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h6c: begin
							r_fld_res_9_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_err_10 <= w_sys_tmp1;

									end
								end

							endcase
						end

						7'h5f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_err_10 <= w_sys_tmp513;

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h12)) begin
										r_threadTop_err_10 <= w_sys_tmp516;

									end
								end

							endcase
						end

						7'h66: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_threadTop_err_10 <= w_sys_tmp526;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h19: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_alpha_11 <= w_sys_tmp144;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h52: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_sum_12 <= w_sys_tmp404;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b)) begin
										r_threadTop_sum_12 <= w_sys_tmp407;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h33)) begin
										r_threadTop_delta_13 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_threadTop_step==7'h23) || (r_sys_threadTop_step==7'h2b)) begin
										r_threadTop_delta_13 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_threadTop_step==7'h1b) || (r_sys_threadTop_step==7'h1e)) begin
										r_threadTop_delta_13 <= w_sys_tmp309;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h27)) begin
										r_threadTop_delta_13 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_threadTop_step==7'h17) || (r_sys_threadTop_step==7'h19)) begin
										r_threadTop_delta_13 <= w_sys_tmp421;

									end
									else
									if((r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h2f)) begin
										r_threadTop_delta_13 <= r_sys_tmp0_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_i_14 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_i_14 <= w_sys_tmp35;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h9: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_15 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'hf<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h13)) begin
										r_threadTop_j_15 <= w_sys_tmp49;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hf: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_i_16 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h11: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_i_16 <= w_sys_tmp95;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h14: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_17 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'hf<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h13)) begin
										r_threadTop_j_17 <= w_sys_tmp107;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_i_18 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h66: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_i_18 <= w_sys_tmp528;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_19 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_threadTop_j_19 <= w_sys_tmp156;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_20 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h34: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_threadTop_k_20 <= w_sys_tmp249;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_21 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_j_21 <= w_sys_tmp200;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h36: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_22 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_threadTop_k_22 <= w_sys_tmp304;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h3c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_23 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_j_23 <= w_sys_tmp263;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h43: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_24 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_24 <= w_sys_tmp306;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h48: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_25 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_j_25 <= w_sys_tmp328;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_l_26 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h50: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_l_26 <= w_sys_tmp403;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h54: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_27 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_threadTop_k_27 <= w_sys_tmp418;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h5a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_28 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_j_28 <= w_sys_tmp439;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h61: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_29 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1)) begin
										r_threadTop_k_29 <= w_sys_tmp525;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy0_j_31 <= r_threadTop_j_19;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_copy0_j_31 <= w_sys_tmp155;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2f: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy0_j_32 <= r_threadTop_j_21;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_copy0_j_32 <= w_sys_tmp199;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h3c: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy0_j_33 <= r_threadTop_j_23;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_copy0_j_33 <= w_sys_tmp262;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h48: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy0_j_34 <= r_threadTop_j_25;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h21) || (r_sys_threadTop_step==7'h29) || (r_sys_threadTop_step==7'h31) || (r_sys_threadTop_step==7'h39)) begin
										r_threadTop_copy0_j_34 <= w_sys_tmp326;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h48: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy1_j_35 <= r_threadTop_j_25;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h20) || (r_sys_threadTop_step==7'h28) || (r_sys_threadTop_step==7'h30) || (r_sys_threadTop_step==7'h38) || (r_sys_threadTop_step==7'h40)) begin
										r_threadTop_copy1_j_35 <= w_sys_tmp327;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h5a: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy0_j_36 <= r_threadTop_j_28;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h25) || (r_sys_threadTop_step==7'h2d) || (r_sys_threadTop_step==7'h35)) begin
										r_threadTop_copy0_j_36 <= w_sys_tmp437;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h5a: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy1_j_37 <= r_threadTop_j_28;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c) || (r_sys_threadTop_step==7'h34) || (r_sys_threadTop_step==7'h3c)) begin
										r_threadTop_copy1_j_37 <= w_sys_tmp438;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp0_float <= w_ip_rand_result_1;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp0_float <= w_ip_rand_result_6;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'ha)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'ha)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_tmp0_float <= w_fld_res_9_dataout_1;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8) || (r_sys_threadTop_step==7'ha)) begin
										r_sys_tmp0_float <= w_fld_hidden_6_dataout_1;

									end
									else
									if((r_sys_threadTop_step==7'h7) || (r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hb) || (r_sys_threadTop_step==7'h1b) || (r_sys_threadTop_step==7'h1f)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp1_float <= w_ip_rand_result_2;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp1_float <= w_ip_rand_result_7;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h9)) begin
										r_sys_tmp1_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h9)) begin
										r_sys_tmp1_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_tmp1_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp2_float <= w_ip_rand_result_4;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp2_float <= w_ip_rand_result_9;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_sys_tmp2_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_sys_tmp2_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_sys_tmp2_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp3_float <= w_ip_rand_result_3;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp3_float <= w_ip_rand_result_8;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp3_float <= w_fld_hidden_6_dataout_1;

									end
									else
									if((r_sys_threadTop_step==7'hb)) begin
										r_sys_tmp3_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h40: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp3_float <= w_fld_output_7_dataout_1;

									end
									else
									if((r_sys_threadTop_step==7'hb)) begin
										r_sys_tmp3_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h4)) begin
										r_sys_tmp3_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp4_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp4_float <= w_fld_output_7_dataout_1;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h4)) begin
										r_sys_tmp4_float <= w_fld_input_5_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp5_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

						7'h58: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h9)) begin
										r_sys_tmp5_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp5_float <= w_fld_w2_4_dataout_1;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp5_float <= w_fld_w1_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp6_float <= w_fld_w2_4_dataout_1;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_sys_tmp6_float <= w_fld_input_5_dataout_1;

									end
								end

							endcase
						end

						7'h65: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7)) begin
										r_sys_tmp6_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6) || (r_sys_threadTop_step==7'hc)) begin
										r_sys_tmp7_float <= w_fld_output_7_dataout_1;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp7_float <= w_fld_input_5_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3) || (r_sys_threadTop_step==7'h5)) begin
										r_sys_tmp8_float <= w_fld_res_9_dataout_1;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp8_float <= w_fld_input_5_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3) || (r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hf)) begin
										r_sys_tmp9_float <= w_fld_output_7_dataout_1;

									end
									else
									if((r_sys_threadTop_step==7'h27)) begin
										r_sys_tmp9_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h5e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_tmp9_float <= w_fld_input_5_dataout_1;

									end
									else
									if((r_sys_threadTop_step==7'h1d)) begin
										r_sys_tmp9_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'hf) || (r_sys_threadTop_step==7'h12) || (r_sys_threadTop_step==7'h15)) begin
										r_sys_tmp10_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_sys_tmp10_float <= w_fld_res_9_dataout_1;

									end
									else
									if((r_sys_threadTop_step==7'h21) || (r_sys_threadTop_step==7'h24)) begin
										r_sys_tmp10_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
