/*
TimeStamp:	2016/9/9		16:52
*/


module subunder(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	input  signed  [14:0] i_fld_u_0_addr_0,	
	input          [31:0] i_fld_u_0_datain_0,	
	output         [31:0] o_fld_u_0_dataout_0,	
	input                 i_fld_u_0_r_w_0,	
	input  signed  [14:0] i_fld_result_1_addr_0,	
	input          [31:0] i_fld_result_1_datain_0,	
	output         [31:0] o_fld_result_1_dataout_0,	
	input                 i_fld_result_1_r_w_0	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 3:0] r_sys_run_phase;
	reg         [ 1:0] r_sys_run_stage;
	reg         [ 7:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 1:0] w_sys_run_stage_p1;
	wire        [ 7:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	wire signed [14:0] w_fld_result_1_addr_0;
	wire        [31:0] w_fld_result_1_datain_0;
	wire        [31:0] w_fld_result_1_dataout_0;
	wire               w_fld_result_1_r_w_0;
	wire               w_fld_result_1_ce_0;
	reg  signed [14:0] r_fld_result_1_addr_1;
	reg         [31:0] r_fld_result_1_datain_1;
	wire        [31:0] w_fld_result_1_dataout_1;
	reg                r_fld_result_1_r_w_1;
	wire               w_fld_result_1_ce_1;
	reg         [31:0] r_fld_r1_2;
	reg         [31:0] r_fld_r2_3;
	reg         [31:0] r_fld_dx_4;
	reg         [31:0] r_fld_dy_5;
	reg         [31:0] r_fld_dt_6;
	reg  signed [31:0] r_run_k_7;
	reg  signed [31:0] r_run_j_8;
	reg  signed [31:0] r_run_copy0_j_9;
	reg  signed [31:0] r_run_copy1_j_10;
	reg  signed [31:0] r_run_copy2_j_11;
	reg  signed [31:0] r_run_copy3_j_12;
	reg  signed [31:0] r_run_copy4_j_13;
	reg  signed [31:0] r_run_copy5_j_14;
	reg  signed [31:0] r_run_copy6_j_15;
	reg  signed [31:0] r_run_copy7_j_16;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	reg         [31:0] r_sys_tmp48_float;
	reg         [31:0] r_sys_tmp49_float;
	reg         [31:0] r_sys_tmp50_float;
	reg         [31:0] r_sys_tmp51_float;
	reg         [31:0] r_sys_tmp52_float;
	reg         [31:0] r_sys_tmp53_float;
	reg         [31:0] r_sys_tmp54_float;
	reg         [31:0] r_sys_tmp55_float;
	reg         [31:0] r_sys_tmp56_float;
	reg         [31:0] r_sys_tmp57_float;
	reg         [31:0] r_sys_tmp58_float;
	reg         [31:0] r_sys_tmp59_float;
	reg         [31:0] r_sys_tmp60_float;
	reg         [31:0] r_sys_tmp61_float;
	reg         [31:0] r_sys_tmp62_float;
	reg         [31:0] r_sys_tmp63_float;
	reg         [31:0] r_sys_tmp64_float;
	reg         [31:0] r_sys_tmp65_float;
	reg         [31:0] r_sys_tmp66_float;
	reg         [31:0] r_sys_tmp67_float;
	reg         [31:0] r_sys_tmp68_float;
	reg         [31:0] r_sys_tmp69_float;
	reg         [31:0] r_sys_tmp70_float;
	reg         [31:0] r_sys_tmp71_float;
	reg         [31:0] r_sys_tmp72_float;
	wire        [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp4;
	wire signed [31:0] w_sys_tmp6;
	wire               w_sys_tmp7;
	wire               w_sys_tmp8;
	wire signed [31:0] w_sys_tmp9;
	wire signed [31:0] w_sys_tmp10;
	wire signed [31:0] w_sys_tmp11;
	wire               w_sys_tmp12;
	wire               w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire signed [31:0] w_sys_tmp17;
	wire signed [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire        [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire signed [31:0] w_sys_tmp22;
	wire        [31:0] w_sys_tmp24;
	wire signed [31:0] w_sys_tmp26;
	wire signed [31:0] w_sys_tmp27;
	wire signed [31:0] w_sys_tmp28;
	wire        [31:0] w_sys_tmp31;
	wire        [31:0] w_sys_tmp32;
	wire signed [31:0] w_sys_tmp33;
	wire signed [31:0] w_sys_tmp34;
	wire signed [31:0] w_sys_tmp36;
	wire signed [31:0] w_sys_tmp37;
	wire signed [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp43;
	wire signed [31:0] w_sys_tmp44;
	wire signed [31:0] w_sys_tmp49;
	wire signed [31:0] w_sys_tmp50;
	wire signed [31:0] w_sys_tmp52;
	wire signed [31:0] w_sys_tmp53;
	wire signed [31:0] w_sys_tmp54;
	wire        [31:0] w_sys_tmp56;
	wire signed [31:0] w_sys_tmp57;
	wire signed [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp59;
	wire signed [31:0] w_sys_tmp60;
	wire signed [31:0] w_sys_tmp61;
	wire signed [31:0] w_sys_tmp62;
	wire signed [31:0] w_sys_tmp63;
	wire signed [31:0] w_sys_tmp64;
	wire signed [31:0] w_sys_tmp66;
	wire signed [31:0] w_sys_tmp67;
	wire        [31:0] w_sys_tmp1057;
	wire        [31:0] w_sys_tmp1058;
	wire        [31:0] w_sys_tmp1059;
	wire        [31:0] w_sys_tmp1060;
	wire        [31:0] w_sys_tmp1061;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 2'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 8'h1);
	assign o_fld_u_0_dataout_0 = w_fld_u_0_dataout_0;
	assign w_fld_u_0_addr_0 = i_fld_u_0_addr_0;
	assign w_fld_u_0_datain_0 = i_fld_u_0_datain_0;
	assign w_fld_u_0_r_w_0 = i_fld_u_0_r_w_0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign o_fld_result_1_dataout_0 = w_fld_result_1_dataout_0;
	assign w_fld_result_1_addr_0 = i_fld_result_1_addr_0;
	assign w_fld_result_1_datain_0 = i_fld_result_1_datain_0;
	assign w_fld_result_1_r_w_0 = i_fld_result_1_r_w_0;
	assign w_fld_result_1_ce_0 = w_sys_ce;
	assign w_fld_result_1_ce_1 = w_sys_ce;
	assign w_sys_tmp1 = 32'h3c000000;
	assign w_sys_tmp3 = 32'h3ba3d70a;
	assign w_sys_tmp4 = 32'h42a3d70a;
	assign w_sys_tmp6 = 32'sh00000041;
	assign w_sys_tmp7 = ( !w_sys_tmp8 );
	assign w_sys_tmp8 = (w_sys_tmp9 < r_run_k_7);
	assign w_sys_tmp9 = 32'sh00000080;
	assign w_sys_tmp10 = (r_run_k_7 + w_sys_intOne);
	assign w_sys_tmp11 = 32'sh00000002;
	assign w_sys_tmp12 = ( !w_sys_tmp13 );
	assign w_sys_tmp13 = (w_sys_tmp14 < r_run_j_8);
	assign w_sys_tmp14 = 32'sh00000080;
	assign w_sys_tmp17 = (w_sys_tmp18 + r_run_k_7);
	assign w_sys_tmp18 = (r_run_j_8 * w_sys_tmp19);
	assign w_sys_tmp19 = 32'sh00000081;
	assign w_sys_tmp20 = w_ip_AddFloat_result_0;
	assign w_sys_tmp21 = (w_sys_tmp22 + r_run_k_7);
	assign w_sys_tmp22 = (r_run_copy7_j_16 * w_sys_tmp19);
	assign w_sys_tmp24 = w_ip_MultFloat_product_0;
	assign w_sys_tmp26 = (w_sys_tmp27 + r_run_k_7);
	assign w_sys_tmp27 = (w_sys_tmp28 * w_sys_tmp19);
	assign w_sys_tmp28 = (r_run_copy6_j_15 + w_sys_intOne);
	assign w_sys_tmp31 = 32'h40000000;
	assign w_sys_tmp32 = w_fld_u_0_dataout_1;
	assign w_sys_tmp33 = (w_sys_tmp34 + r_run_k_7);
	assign w_sys_tmp34 = (r_run_copy5_j_14 * w_sys_tmp19);
	assign w_sys_tmp36 = (w_sys_tmp37 + r_run_k_7);
	assign w_sys_tmp37 = (w_sys_tmp38 * w_sys_tmp19);
	assign w_sys_tmp38 = (r_run_copy4_j_13 - w_sys_intOne);
	assign w_sys_tmp42 = (w_sys_tmp43 + w_sys_intOne);
	assign w_sys_tmp43 = (w_sys_tmp44 + r_run_k_7);
	assign w_sys_tmp44 = (r_run_copy3_j_12 * w_sys_tmp19);
	assign w_sys_tmp49 = (w_sys_tmp50 + r_run_k_7);
	assign w_sys_tmp50 = (r_run_copy2_j_11 * w_sys_tmp19);
	assign w_sys_tmp52 = (w_sys_tmp53 - w_sys_intOne);
	assign w_sys_tmp53 = (w_sys_tmp54 + r_run_k_7);
	assign w_sys_tmp54 = (r_run_copy1_j_10 * w_sys_tmp19);
	assign w_sys_tmp56 = 32'h42c80000;
	assign w_sys_tmp57 = (r_run_copy0_j_9 - w_sys_intOne);
	assign w_sys_tmp58 = (r_run_k_7 - w_sys_intOne);
	assign w_sys_tmp59 = (r_run_copy0_j_9 + w_sys_intOne);
	assign w_sys_tmp60 = (r_run_copy1_j_10 + w_sys_intOne);
	assign w_sys_tmp61 = (r_run_copy2_j_11 + w_sys_intOne);
	assign w_sys_tmp62 = (r_run_copy3_j_12 + w_sys_intOne);
	assign w_sys_tmp63 = (r_run_copy4_j_13 + w_sys_intOne);
	assign w_sys_tmp64 = (r_run_copy5_j_14 + w_sys_intOne);
	assign w_sys_tmp66 = (r_run_copy7_j_16 + w_sys_intOne);
	assign w_sys_tmp67 = (r_run_j_8 + w_sys_intOne);
	assign w_sys_tmp1057 = 32'h0;
	assign w_sys_tmp1058 = 32'h0;
	assign w_sys_tmp1059 = 32'h0;
	assign w_sys_tmp1060 = 32'h0;
	assign w_sys_tmp1061 = 32'h0;


	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_result_1(
			.clk (clock),
			.ce_0 (w_fld_result_1_ce_0),
			.addr_0 (w_fld_result_1_addr_0),
			.datain_0 (w_fld_result_1_datain_0),
			.dataout_0 (w_fld_result_1_dataout_0),
			.r_w_0 (w_fld_result_1_r_w_0),
			.ce_1 (w_fld_result_1_ce_1),
			.addr_1 (r_fld_result_1_addr_1),
			.datain_1 (r_fld_result_1_datain_1),
			.dataout_1 (w_fld_result_1_dataout_1),
			.r_w_1 (r_fld_result_1_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h21) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h67)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==8'h51) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'ha3)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==8'h37) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'hb4)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==8'h76) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'had)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h96)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp20;

									end
									else
									if((r_sys_run_step==8'h7c) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h91)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==8'h71) || (r_sys_run_step==8'hab)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==8'h5c) || (r_sys_run_step==8'hae)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==8'h1e) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h8e)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==8'h6d) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'haa)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==8'h1d) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h89)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==8'ha7)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==8'h47) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'hb3)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==8'h7f) || (r_sys_run_step==8'hb0) || (r_sys_run_step==8'hb6) || (r_sys_run_step==8'hb8)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==8'h8d)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h95)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==8'h1a) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h9f)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==8'h63) || (r_sys_run_step==8'ha0)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h9a)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==8'h66) || (r_sys_run_step==8'h92)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==8'h6a) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'hb1) || (r_sys_run_step==8'hb7)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==8'h7b) || (r_sys_run_step==8'h9e)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h82)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==8'h40) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'hb5)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==8'h10) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h90)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==8'hc) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'ha4)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp70_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h88)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==8'h8a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h89) || (r_sys_run_step==8'h8b)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h23) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h73)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h11) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h77)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==8'h1d) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'h94) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'h9f) || (r_sys_run_step==8'ha0) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'ha4) || (r_sys_run_step==8'ha5) || (r_sys_run_step==8'ha7) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'haa) || (r_sys_run_step==8'hab) || (r_sys_run_step==8'had) || (r_sys_run_step==8'hae) || (r_sys_run_step==8'hb0) || (r_sys_run_step==8'hb1) || (8'hb3<=r_sys_run_step && r_sys_run_step<=8'hb8)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp24;

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h8e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h15) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h81)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h70) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h8f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h5c) || (r_sys_run_step==8'h63)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==8'h91)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h90) || (r_sys_run_step==8'h92)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==8'h26) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h93)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==8'h40) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h68)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h35) || (r_sys_run_step==8'h84)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h1c) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h6c)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h2d) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'h96)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h7f) || (r_sys_run_step==8'h82)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h4d) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h65)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==8'h78) || (r_sys_run_step==8'h7b)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==8'h97)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp24[31], w_sys_tmp24[30:0] };

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp50_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'had) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hb3)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==8'h1b) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'hab)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==8'h67) || (r_sys_run_step==8'h8e)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==8'h47) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h94)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h55) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h9e)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==8'h32) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'ha0) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'ha6) || (r_sys_run_step==8'ha9) || (r_sys_run_step==8'hac)) begin
										r_ip_MultFloat_multiplicand_0 <= r_fld_r2_3;

									end
									else
									if((r_sys_run_step==8'h4) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8c)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp31;

									end
									else
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'ha7) || (r_sys_run_step==8'hb1)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==8'h33) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h9c)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==8'h57) || (r_sys_run_step==8'h7f)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==8'h4e) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h99)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'ha4) || (r_sys_run_step==8'haf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==8'h36) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h86)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==8'hd) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'hb0)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h8d)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp48_float;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h52)) begin
										r_ip_MultFloat_multiplicand_0 <= r_fld_dt_6;

									end
									else
									if((r_sys_run_step==8'h28) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'haa)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'h9f)) begin
										r_ip_MultFloat_multiplicand_0 <= r_fld_r1_2;

									end
									else
									if((r_sys_run_step==8'h22) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'ha5)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==8'h1d) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'ha2) || (r_sys_run_step==8'hae)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp51_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hb3)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h99)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==8'h17) || (r_sys_run_step==8'h79)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp20;

									end
									else
									if((r_sys_run_step==8'h92)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'h9c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h45) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h9f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==8'h1d) || (r_sys_run_step==8'h8f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp31_float;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h52)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp56;

									end
									else
									if((r_sys_run_step==8'h2d) || (r_sys_run_step==8'hb2)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==8'h3a) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'ha3)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==8'haf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'ha8)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h7d)) begin
										r_ip_MultFloat_multiplier_0 <= r_fld_dx_4;

									end
									else
									if((r_sys_run_step==8'h4e) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h90)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==8'h6c) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h95)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==8'h32) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'ha0)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==8'h8d)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==8'h18) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h9a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==8'hb0)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'ha5)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h36) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h8e) || (r_sys_run_step==8'h93) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'h9d) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'ha4) || (r_sys_run_step==8'ha7) || (r_sys_run_step==8'haa) || (r_sys_run_step==8'had)) begin
										r_ip_MultFloat_multiplier_0 <= r_fld_dy_5;

									end
									else
									if((r_sys_run_step==8'h59) || (r_sys_run_step==8'h61)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==8'h28) || (r_sys_run_step==8'hab)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==8'h5d) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'ha6)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==8'h9b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==8'h22) || (r_sys_run_step==8'h97)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'hb1)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h8b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==8'ha2)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h94)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'h34) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'ha9)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==8'h4) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8c)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp32;

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h29) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'hac)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'h9e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'hae)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp14_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h1c) || (8'h1e<=r_sys_run_step && r_sys_run_step<=8'h27)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp58;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp57;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						4'hf: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h0: begin
							r_sys_run_phase <= 4'h2;
						end

						4'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 4'h4;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 4'h5;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7) ? 4'h9 : 4'hf);

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 4'h5;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 4'ha;

									end
								end

							endcase
						end

						4'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12) ? 4'hd : 4'h6);

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hbd)) begin
										r_sys_run_phase <= 4'ha;

									end
								end

							endcase
						end

						4'hf: begin
							r_sys_run_phase <= 4'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						4'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hbd)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 8'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						4'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						4'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						4'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						4'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'hbc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'hbd)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						4'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						4'hf: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h88)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp36[14:0] );

									end
									else
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp52[14:0] );

									end
									else
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h8a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp49[14:0] );

									end
									else
									if((r_sys_run_step==8'h4) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h89)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp42[14:0] );

									end
									else
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h87)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp33[14:0] );

									end
									else
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h86)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp26[14:0] );

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h85)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp21[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h8b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						4'hf: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_result_1_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6b) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'haf) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hb5) || (8'hb8<=r_sys_run_step && r_sys_run_step<=8'hbd)) begin
										r_fld_result_1_addr_1 <= $signed( w_sys_tmp17[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6b) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'haf) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hb5) || (8'hb8<=r_sys_run_step && r_sys_run_step<=8'hbd)) begin
										r_fld_result_1_datain_1 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_result_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6b) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'haf) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hb5) || (8'hb8<=r_sys_run_step && r_sys_run_step<=8'hbd)) begin
										r_fld_result_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						4'hf: begin
							r_fld_result_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_r1_2 <= w_sys_tmp1057;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_r1_2 <= w_sys_tmp4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_r2_3 <= w_sys_tmp1058;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_r2_3 <= w_sys_tmp4;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_dx_4 <= w_sys_tmp1059;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_dx_4 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_dy_5 <= w_sys_tmp1060;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_dy_5 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_dt_6 <= w_sys_tmp1061;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_dt_6 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_7 <= w_sys_tmp6;

									end
								end

							endcase
						end

						4'h6: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_7 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h9: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_8 <= w_sys_tmp11;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6b) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'h99) || (r_sys_run_step==8'h9e) || (r_sys_run_step==8'ha3) || (r_sys_run_step==8'ha8) || (r_sys_run_step==8'hac) || (r_sys_run_step==8'haf) || (r_sys_run_step==8'hb2) || (r_sys_run_step==8'hb5) || (8'hb8<=r_sys_run_step && r_sys_run_step<=8'hbd)) begin
										r_run_j_8 <= w_sys_tmp67;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_9 <= r_run_j_8;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h1d)) begin
										r_run_copy0_j_9 <= w_sys_tmp59;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy1_j_10 <= r_run_j_8;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8b)) begin
										r_run_copy1_j_10 <= w_sys_tmp60;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy2_j_11 <= r_run_j_8;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h8a)) begin
										r_run_copy2_j_11 <= w_sys_tmp61;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy3_j_12 <= r_run_j_8;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h4) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h20) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h89)) begin
										r_run_copy3_j_12 <= w_sys_tmp62;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy4_j_13 <= r_run_j_8;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h88)) begin
										r_run_copy4_j_13 <= w_sys_tmp63;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy5_j_14 <= r_run_j_8;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h87)) begin
										r_run_copy5_j_14 <= w_sys_tmp64;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy6_j_15 <= r_run_j_8;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h86)) begin
										r_run_copy6_j_15 <= w_sys_tmp28;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'h9: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy7_j_16 <= r_run_j_8;

									end
								end

							endcase
						end

						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h1c) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h85)) begin
										r_run_copy7_j_16 <= w_sys_tmp66;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2e)) begin
										r_sys_tmp0_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2c)) begin
										r_sys_tmp1_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2b)) begin
										r_sys_tmp2_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2a)) begin
										r_sys_tmp3_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h29)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h27)) begin
										r_sys_tmp5_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h26)) begin
										r_sys_tmp6_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h25)) begin
										r_sys_tmp7_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h24)) begin
										r_sys_tmp8_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h23)) begin
										r_sys_tmp9_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h21)) begin
										r_sys_tmp10_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_tmp11_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1f)) begin
										r_sys_tmp12_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_tmp13_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1c)) begin
										r_sys_tmp14_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sys_tmp15_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sys_tmp16_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_sys_tmp17_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sys_tmp18_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp19_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sys_tmp20_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h13)) begin
										r_sys_tmp21_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_tmp22_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h11)) begin
										r_sys_tmp23_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5a) || (r_sys_run_step==8'h80)) begin
										r_sys_tmp24_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h55) || (r_sys_run_step==8'h7d)) begin
										r_sys_tmp25_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h4d) || (r_sys_run_step==8'h54)) begin
										r_sys_tmp26_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h32) || (r_sys_run_step==8'h58)) begin
										r_sys_tmp27_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hb) || (r_sys_run_step==8'h2d)) begin
										r_sys_tmp28_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'h28)) begin
										r_sys_tmp29_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h9) || (r_sys_run_step==8'h22)) begin
										r_sys_tmp30_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'h1d)) begin
										r_sys_tmp31_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'h17)) begin
										r_sys_tmp32_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h43)) begin
										r_sys_tmp33_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_sys_tmp33_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_tmp34_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_sys_tmp34_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h45) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h97)) begin
										r_sys_tmp35_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h42) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6a)) begin
										r_sys_tmp36_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2b) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h7d)) begin
										r_sys_tmp37_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h27) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h74)) begin
										r_sys_tmp38_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2b) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h9c)) begin
										r_sys_tmp39_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1c) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h5f)) begin
										r_sys_tmp40_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h19) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h82)) begin
										r_sys_tmp41_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h33) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h89)) begin
										r_sys_tmp42_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h31) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h85)) begin
										r_sys_tmp43_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1d) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h86) || (r_sys_run_step==8'ha4)) begin
										r_sys_tmp44_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hf)) begin
										r_sys_tmp45_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==8'h4e) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h90)) begin
										r_sys_tmp45_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_tmp46_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==8'h3d) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h8e)) begin
										r_sys_tmp46_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h22) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h8d) || (r_sys_run_step==8'haa)) begin
										r_sys_tmp47_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h20) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h68)) begin
										r_sys_tmp48_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h15) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h96) || (r_sys_run_step==8'h9c)) begin
										r_sys_tmp49_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h12) || (r_sys_run_step==8'h23) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h93)) begin
										r_sys_tmp50_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hf) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h8c) || (r_sys_run_step==8'ha2)) begin
										r_sys_tmp51_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'he)) begin
										r_sys_tmp52_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==8'h4b) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'h9f)) begin
										r_sys_tmp52_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_sys_tmp53_float <= w_ip_FixedToFloat_floating_0;

									end
									else
									if((r_sys_run_step==8'h36) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h94)) begin
										r_sys_tmp53_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2e) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h8a) || (r_sys_run_step==8'h95) || (r_sys_run_step==8'ha5)) begin
										r_sys_tmp54_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h28) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h87) || (r_sys_run_step==8'h9b) || (r_sys_run_step==8'had)) begin
										r_sys_tmp55_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h16) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'ha0) || (r_sys_run_step==8'hb0) || (r_sys_run_step==8'hb6)) begin
										r_sys_tmp56_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hb) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h97) || (r_sys_run_step==8'hac)) begin
										r_sys_tmp57_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5b) || (r_sys_run_step==8'h62)) begin
										r_sys_tmp58_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==8'h76) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h8b)) begin
										r_sys_tmp58_float <= w_fld_u_0_dataout_1;

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sys_tmp58_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'he) || (r_sys_run_step==8'h1b) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h9d)) begin
										r_sys_tmp59_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h1b) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h86)) begin
										r_sys_tmp60_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'hd) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h72)) begin
										r_sys_tmp61_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h8) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h79)) begin
										r_sys_tmp62_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h7) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h98) || (r_sys_run_step==8'ha9)) begin
										r_sys_tmp63_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h8f) || (r_sys_run_step==8'h90) || (r_sys_run_step==8'h92) || (r_sys_run_step==8'ha6)) begin
										r_sys_tmp64_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h8d)) begin
										r_sys_tmp65_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h1d) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h8a)) begin
										r_sys_tmp66_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h14) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h80)) begin
										r_sys_tmp67_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h13) || (r_sys_run_step==8'h1a) || (r_sys_run_step==8'h21) || (r_sys_run_step==8'h24) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h91) || (r_sys_run_step==8'h9a) || (r_sys_run_step==8'ha9) || (r_sys_run_step==8'hb3)) begin
										r_sys_tmp68_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'ha) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h6b)) begin
										r_sys_tmp69_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h6) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1f) || (r_sys_run_step==8'h25) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h87)) begin
										r_sys_tmp70_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h22) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h88) || (r_sys_run_step==8'h89) || (r_sys_run_step==8'h8b) || (r_sys_run_step==8'ha1) || (r_sys_run_step==8'haf) || (r_sys_run_step==8'hb2)) begin
										r_sys_tmp71_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						4'hd: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==8'h5) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h18) || (r_sys_run_step==8'h1e) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h88)) begin
										r_sys_tmp72_float <= w_fld_u_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
