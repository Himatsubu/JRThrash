/*
TimeStamp:	2016/9/12		16:35
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	output signed  [31:0] o_run_return	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [31:0] r_sys_run_return;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 5:0] r_sys_run_phase;
	reg         [ 3:0] r_sys_run_stage;
	reg         [ 7:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 3:0] w_sys_run_stage_p1;
	wire        [ 7:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_9;
	reg  signed [31:0] r_run_j_10;
	reg  signed [31:0] r_run_n_11;
	reg  signed [31:0] r_run_mx_12;
	reg  signed [31:0] r_run_my_13;
	reg  signed [31:0] r_run_nlast_14;
	reg         [31:0] r_run_dx_15;
	reg         [31:0] r_run_dy_16;
	reg         [31:0] r_run_dt_17;
	reg         [31:0] r_run_r1_18;
	reg         [31:0] r_run_r2_19;
	reg  signed [31:0] r_run_copy0_j_20;
	reg  signed [31:0] r_run_copy1_j_21;
	reg  signed [31:0] r_run_copy2_j_22;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [14:0] w_sub03_u_addr;
	reg  signed [14:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [14:0] w_sub03_result_addr;
	reg  signed [14:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [14:0] w_sub02_u_addr;
	reg  signed [14:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [14:0] w_sub02_result_addr;
	reg  signed [14:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [14:0] w_sub01_u_addr;
	reg  signed [14:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [14:0] w_sub01_result_addr;
	reg  signed [14:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [14:0] w_sub00_u_addr;
	reg  signed [14:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [14:0] w_sub00_result_addr;
	reg  signed [14:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [14:0] w_sub07_u_addr;
	reg  signed [14:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [14:0] w_sub07_result_addr;
	reg  signed [14:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [14:0] w_sub06_u_addr;
	reg  signed [14:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [14:0] w_sub06_result_addr;
	reg  signed [14:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [14:0] w_sub05_u_addr;
	reg  signed [14:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [14:0] w_sub05_result_addr;
	reg  signed [14:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [14:0] w_sub04_u_addr;
	reg  signed [14:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [14:0] w_sub04_result_addr;
	reg  signed [14:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	reg         [31:0] r_sys_tmp48_float;
	reg         [31:0] r_sys_tmp49_float;
	reg         [31:0] r_sys_tmp50_float;
	reg         [31:0] r_sys_tmp51_float;
	reg         [31:0] r_sys_tmp52_float;
	reg         [31:0] r_sys_tmp53_float;
	reg         [31:0] r_sys_tmp54_float;
	reg         [31:0] r_sys_tmp55_float;
	reg         [31:0] r_sys_tmp56_float;
	reg         [31:0] r_sys_tmp57_float;
	reg         [31:0] r_sys_tmp58_float;
	reg         [31:0] r_sys_tmp59_float;
	reg         [31:0] r_sys_tmp60_float;
	reg         [31:0] r_sys_tmp61_float;
	reg         [31:0] r_sys_tmp62_float;
	reg         [31:0] r_sys_tmp63_float;
	reg         [31:0] r_sys_tmp64_float;
	reg         [31:0] r_sys_tmp65_float;
	reg         [31:0] r_sys_tmp66_float;
	reg         [31:0] r_sys_tmp67_float;
	reg         [31:0] r_sys_tmp68_float;
	reg         [31:0] r_sys_tmp69_float;
	reg         [31:0] r_sys_tmp70_float;
	reg         [31:0] r_sys_tmp71_float;
	reg         [31:0] r_sys_tmp72_float;
	reg         [31:0] r_sys_tmp73_float;
	reg         [31:0] r_sys_tmp74_float;
	reg         [31:0] r_sys_tmp75_float;
	reg         [31:0] r_sys_tmp76_float;
	reg         [31:0] r_sys_tmp77_float;
	reg         [31:0] r_sys_tmp78_float;
	reg         [31:0] r_sys_tmp79_float;
	reg         [31:0] r_sys_tmp80_float;
	reg         [31:0] r_sys_tmp81_float;
	reg         [31:0] r_sys_tmp82_float;
	reg         [31:0] r_sys_tmp83_float;
	reg         [31:0] r_sys_tmp84_float;
	reg         [31:0] r_sys_tmp85_float;
	reg         [31:0] r_sys_tmp86_float;
	reg         [31:0] r_sys_tmp87_float;
	reg         [31:0] r_sys_tmp88_float;
	reg         [31:0] r_sys_tmp89_float;
	reg         [31:0] r_sys_tmp90_float;
	reg         [31:0] r_sys_tmp91_float;
	reg         [31:0] r_sys_tmp92_float;
	reg         [31:0] r_sys_tmp93_float;
	reg         [31:0] r_sys_tmp94_float;
	wire signed [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire               w_sys_tmp8;
	wire               w_sys_tmp9;
	wire signed [31:0] w_sys_tmp10;
	wire               w_sys_tmp11;
	wire               w_sys_tmp12;
	wire signed [31:0] w_sys_tmp15;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire        [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp19;
	wire               w_sys_tmp56;
	wire               w_sys_tmp57;
	wire signed [31:0] w_sys_tmp58;
	wire               w_sys_tmp59;
	wire               w_sys_tmp60;
	wire signed [31:0] w_sys_tmp63;
	wire signed [31:0] w_sys_tmp64;
	wire        [31:0] w_sys_tmp65;
	wire signed [31:0] w_sys_tmp67;
	wire signed [31:0] w_sys_tmp68;
	wire        [31:0] w_sys_tmp70;
	wire signed [31:0] w_sys_tmp72;
	wire signed [31:0] w_sys_tmp73;
	wire        [31:0] w_sys_tmp75;
	wire signed [31:0] w_sys_tmp77;
	wire signed [31:0] w_sys_tmp78;
	wire signed [31:0] w_sys_tmp79;
	wire signed [31:0] w_sys_tmp81;
	wire signed [31:0] w_sys_tmp82;
	wire signed [31:0] w_sys_tmp83;
	wire signed [31:0] w_sys_tmp84;
	wire               w_sys_tmp223;
	wire               w_sys_tmp224;
	wire signed [31:0] w_sys_tmp225;
	wire signed [31:0] w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire        [31:0] w_sys_tmp230;
	wire signed [31:0] w_sys_tmp234;
	wire signed [31:0] w_sys_tmp235;
	wire signed [31:0] w_sys_tmp240;
	wire signed [31:0] w_sys_tmp241;
	wire signed [31:0] w_sys_tmp246;
	wire signed [31:0] w_sys_tmp247;
	wire signed [31:0] w_sys_tmp252;
	wire signed [31:0] w_sys_tmp253;
	wire signed [31:0] w_sys_tmp258;
	wire signed [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp264;
	wire signed [31:0] w_sys_tmp265;
	wire signed [31:0] w_sys_tmp270;
	wire signed [31:0] w_sys_tmp271;
	wire signed [31:0] w_sys_tmp276;
	wire signed [31:0] w_sys_tmp277;
	wire signed [31:0] w_sys_tmp282;
	wire signed [31:0] w_sys_tmp283;
	wire signed [31:0] w_sys_tmp288;
	wire signed [31:0] w_sys_tmp289;
	wire signed [31:0] w_sys_tmp294;
	wire signed [31:0] w_sys_tmp295;
	wire signed [31:0] w_sys_tmp300;
	wire signed [31:0] w_sys_tmp301;
	wire signed [31:0] w_sys_tmp306;
	wire signed [31:0] w_sys_tmp307;
	wire signed [31:0] w_sys_tmp312;
	wire signed [31:0] w_sys_tmp313;
	wire signed [31:0] w_sys_tmp318;
	wire signed [31:0] w_sys_tmp319;
	wire signed [31:0] w_sys_tmp324;
	wire signed [31:0] w_sys_tmp325;
	wire signed [31:0] w_sys_tmp330;
	wire signed [31:0] w_sys_tmp331;
	wire signed [31:0] w_sys_tmp336;
	wire signed [31:0] w_sys_tmp337;
	wire signed [31:0] w_sys_tmp342;
	wire signed [31:0] w_sys_tmp343;
	wire signed [31:0] w_sys_tmp348;
	wire signed [31:0] w_sys_tmp349;
	wire signed [31:0] w_sys_tmp354;
	wire signed [31:0] w_sys_tmp355;
	wire signed [31:0] w_sys_tmp360;
	wire signed [31:0] w_sys_tmp361;
	wire signed [31:0] w_sys_tmp366;
	wire signed [31:0] w_sys_tmp367;
	wire signed [31:0] w_sys_tmp372;
	wire signed [31:0] w_sys_tmp373;
	wire signed [31:0] w_sys_tmp378;
	wire signed [31:0] w_sys_tmp379;
	wire signed [31:0] w_sys_tmp384;
	wire signed [31:0] w_sys_tmp385;
	wire signed [31:0] w_sys_tmp390;
	wire signed [31:0] w_sys_tmp391;
	wire signed [31:0] w_sys_tmp396;
	wire signed [31:0] w_sys_tmp397;
	wire signed [31:0] w_sys_tmp402;
	wire signed [31:0] w_sys_tmp403;
	wire signed [31:0] w_sys_tmp408;
	wire signed [31:0] w_sys_tmp409;
	wire signed [31:0] w_sys_tmp414;
	wire signed [31:0] w_sys_tmp415;
	wire signed [31:0] w_sys_tmp420;
	wire signed [31:0] w_sys_tmp421;
	wire signed [31:0] w_sys_tmp432;
	wire signed [31:0] w_sys_tmp433;
	wire signed [31:0] w_sys_tmp438;
	wire signed [31:0] w_sys_tmp439;
	wire signed [31:0] w_sys_tmp450;
	wire signed [31:0] w_sys_tmp451;
	wire signed [31:0] w_sys_tmp456;
	wire signed [31:0] w_sys_tmp457;
	wire signed [31:0] w_sys_tmp462;
	wire signed [31:0] w_sys_tmp463;
	wire signed [31:0] w_sys_tmp468;
	wire signed [31:0] w_sys_tmp469;
	wire signed [31:0] w_sys_tmp474;
	wire signed [31:0] w_sys_tmp475;
	wire signed [31:0] w_sys_tmp480;
	wire signed [31:0] w_sys_tmp481;
	wire signed [31:0] w_sys_tmp486;
	wire signed [31:0] w_sys_tmp487;
	wire signed [31:0] w_sys_tmp492;
	wire signed [31:0] w_sys_tmp493;
	wire signed [31:0] w_sys_tmp498;
	wire signed [31:0] w_sys_tmp499;
	wire signed [31:0] w_sys_tmp504;
	wire signed [31:0] w_sys_tmp505;
	wire signed [31:0] w_sys_tmp510;
	wire signed [31:0] w_sys_tmp511;
	wire signed [31:0] w_sys_tmp516;
	wire signed [31:0] w_sys_tmp517;
	wire signed [31:0] w_sys_tmp522;
	wire signed [31:0] w_sys_tmp523;
	wire signed [31:0] w_sys_tmp528;
	wire signed [31:0] w_sys_tmp529;
	wire signed [31:0] w_sys_tmp534;
	wire signed [31:0] w_sys_tmp535;
	wire signed [31:0] w_sys_tmp540;
	wire signed [31:0] w_sys_tmp541;
	wire signed [31:0] w_sys_tmp546;
	wire signed [31:0] w_sys_tmp547;
	wire signed [31:0] w_sys_tmp552;
	wire signed [31:0] w_sys_tmp553;
	wire signed [31:0] w_sys_tmp558;
	wire signed [31:0] w_sys_tmp559;
	wire signed [31:0] w_sys_tmp564;
	wire signed [31:0] w_sys_tmp565;
	wire signed [31:0] w_sys_tmp570;
	wire signed [31:0] w_sys_tmp571;
	wire signed [31:0] w_sys_tmp576;
	wire signed [31:0] w_sys_tmp577;
	wire signed [31:0] w_sys_tmp582;
	wire signed [31:0] w_sys_tmp583;
	wire signed [31:0] w_sys_tmp588;
	wire signed [31:0] w_sys_tmp589;
	wire signed [31:0] w_sys_tmp594;
	wire signed [31:0] w_sys_tmp595;
	wire signed [31:0] w_sys_tmp600;
	wire signed [31:0] w_sys_tmp601;
	wire signed [31:0] w_sys_tmp606;
	wire signed [31:0] w_sys_tmp607;
	wire signed [31:0] w_sys_tmp612;
	wire signed [31:0] w_sys_tmp613;
	wire signed [31:0] w_sys_tmp618;
	wire signed [31:0] w_sys_tmp619;
	wire signed [31:0] w_sys_tmp624;
	wire signed [31:0] w_sys_tmp625;
	wire signed [31:0] w_sys_tmp630;
	wire signed [31:0] w_sys_tmp631;
	wire signed [31:0] w_sys_tmp636;
	wire signed [31:0] w_sys_tmp637;
	wire signed [31:0] w_sys_tmp642;
	wire signed [31:0] w_sys_tmp643;
	wire signed [31:0] w_sys_tmp648;
	wire signed [31:0] w_sys_tmp649;
	wire signed [31:0] w_sys_tmp654;
	wire signed [31:0] w_sys_tmp655;
	wire signed [31:0] w_sys_tmp660;
	wire signed [31:0] w_sys_tmp661;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp667;
	wire signed [31:0] w_sys_tmp672;
	wire signed [31:0] w_sys_tmp673;
	wire signed [31:0] w_sys_tmp678;
	wire signed [31:0] w_sys_tmp679;
	wire signed [31:0] w_sys_tmp684;
	wire signed [31:0] w_sys_tmp685;
	wire signed [31:0] w_sys_tmp690;
	wire signed [31:0] w_sys_tmp691;
	wire signed [31:0] w_sys_tmp696;
	wire signed [31:0] w_sys_tmp697;
	wire signed [31:0] w_sys_tmp702;
	wire signed [31:0] w_sys_tmp703;
	wire signed [31:0] w_sys_tmp708;
	wire signed [31:0] w_sys_tmp709;
	wire signed [31:0] w_sys_tmp714;
	wire signed [31:0] w_sys_tmp715;
	wire signed [31:0] w_sys_tmp720;
	wire signed [31:0] w_sys_tmp721;
	wire signed [31:0] w_sys_tmp726;
	wire signed [31:0] w_sys_tmp727;
	wire signed [31:0] w_sys_tmp732;
	wire signed [31:0] w_sys_tmp733;
	wire signed [31:0] w_sys_tmp738;
	wire signed [31:0] w_sys_tmp739;
	wire signed [31:0] w_sys_tmp744;
	wire signed [31:0] w_sys_tmp745;
	wire signed [31:0] w_sys_tmp750;
	wire signed [31:0] w_sys_tmp751;
	wire signed [31:0] w_sys_tmp756;
	wire signed [31:0] w_sys_tmp757;
	wire signed [31:0] w_sys_tmp762;
	wire signed [31:0] w_sys_tmp763;
	wire signed [31:0] w_sys_tmp768;
	wire signed [31:0] w_sys_tmp769;
	wire signed [31:0] w_sys_tmp774;
	wire signed [31:0] w_sys_tmp775;
	wire signed [31:0] w_sys_tmp780;
	wire signed [31:0] w_sys_tmp781;
	wire signed [31:0] w_sys_tmp786;
	wire signed [31:0] w_sys_tmp787;
	wire signed [31:0] w_sys_tmp792;
	wire signed [31:0] w_sys_tmp793;
	wire signed [31:0] w_sys_tmp798;
	wire signed [31:0] w_sys_tmp799;
	wire signed [31:0] w_sys_tmp804;
	wire signed [31:0] w_sys_tmp805;
	wire signed [31:0] w_sys_tmp810;
	wire signed [31:0] w_sys_tmp811;
	wire signed [31:0] w_sys_tmp816;
	wire signed [31:0] w_sys_tmp817;
	wire signed [31:0] w_sys_tmp822;
	wire signed [31:0] w_sys_tmp823;
	wire signed [31:0] w_sys_tmp828;
	wire signed [31:0] w_sys_tmp829;
	wire signed [31:0] w_sys_tmp834;
	wire signed [31:0] w_sys_tmp835;
	wire signed [31:0] w_sys_tmp840;
	wire signed [31:0] w_sys_tmp841;
	wire signed [31:0] w_sys_tmp846;
	wire signed [31:0] w_sys_tmp847;
	wire signed [31:0] w_sys_tmp852;
	wire signed [31:0] w_sys_tmp853;
	wire signed [31:0] w_sys_tmp858;
	wire signed [31:0] w_sys_tmp859;
	wire signed [31:0] w_sys_tmp864;
	wire signed [31:0] w_sys_tmp865;
	wire signed [31:0] w_sys_tmp870;
	wire signed [31:0] w_sys_tmp871;
	wire signed [31:0] w_sys_tmp876;
	wire signed [31:0] w_sys_tmp877;
	wire signed [31:0] w_sys_tmp882;
	wire signed [31:0] w_sys_tmp883;
	wire signed [31:0] w_sys_tmp888;
	wire signed [31:0] w_sys_tmp889;
	wire signed [31:0] w_sys_tmp894;
	wire signed [31:0] w_sys_tmp895;
	wire signed [31:0] w_sys_tmp900;
	wire signed [31:0] w_sys_tmp901;
	wire signed [31:0] w_sys_tmp906;
	wire signed [31:0] w_sys_tmp907;
	wire signed [31:0] w_sys_tmp912;
	wire signed [31:0] w_sys_tmp913;
	wire signed [31:0] w_sys_tmp918;
	wire signed [31:0] w_sys_tmp919;
	wire signed [31:0] w_sys_tmp924;
	wire signed [31:0] w_sys_tmp925;
	wire signed [31:0] w_sys_tmp930;
	wire signed [31:0] w_sys_tmp931;
	wire signed [31:0] w_sys_tmp936;
	wire signed [31:0] w_sys_tmp937;
	wire signed [31:0] w_sys_tmp942;
	wire signed [31:0] w_sys_tmp943;
	wire signed [31:0] w_sys_tmp948;
	wire signed [31:0] w_sys_tmp949;
	wire signed [31:0] w_sys_tmp954;
	wire signed [31:0] w_sys_tmp955;
	wire signed [31:0] w_sys_tmp960;
	wire signed [31:0] w_sys_tmp961;
	wire signed [31:0] w_sys_tmp966;
	wire signed [31:0] w_sys_tmp967;
	wire signed [31:0] w_sys_tmp972;
	wire signed [31:0] w_sys_tmp973;
	wire signed [31:0] w_sys_tmp978;
	wire signed [31:0] w_sys_tmp979;
	wire signed [31:0] w_sys_tmp984;
	wire signed [31:0] w_sys_tmp985;
	wire signed [31:0] w_sys_tmp990;
	wire signed [31:0] w_sys_tmp991;
	wire signed [31:0] w_sys_tmp996;
	wire signed [31:0] w_sys_tmp997;
	wire signed [31:0] w_sys_tmp1002;
	wire signed [31:0] w_sys_tmp1003;
	wire signed [31:0] w_sys_tmp1008;
	wire signed [31:0] w_sys_tmp1009;
	wire signed [31:0] w_sys_tmp1014;
	wire signed [31:0] w_sys_tmp1015;
	wire signed [31:0] w_sys_tmp1020;
	wire signed [31:0] w_sys_tmp1021;
	wire signed [31:0] w_sys_tmp1026;
	wire signed [31:0] w_sys_tmp1027;
	wire signed [31:0] w_sys_tmp1032;
	wire signed [31:0] w_sys_tmp1033;
	wire signed [31:0] w_sys_tmp1037;
	wire signed [31:0] w_sys_tmp1038;
	wire               w_sys_tmp1039;
	wire               w_sys_tmp1040;
	wire signed [31:0] w_sys_tmp1041;
	wire signed [31:0] w_sys_tmp1044;
	wire signed [31:0] w_sys_tmp1045;
	wire        [31:0] w_sys_tmp1046;
	wire signed [31:0] w_sys_tmp1050;
	wire signed [31:0] w_sys_tmp1051;
	wire signed [31:0] w_sys_tmp1056;
	wire signed [31:0] w_sys_tmp1057;
	wire signed [31:0] w_sys_tmp1062;
	wire signed [31:0] w_sys_tmp1063;
	wire signed [31:0] w_sys_tmp1068;
	wire signed [31:0] w_sys_tmp1069;
	wire signed [31:0] w_sys_tmp1074;
	wire signed [31:0] w_sys_tmp1075;
	wire signed [31:0] w_sys_tmp1080;
	wire signed [31:0] w_sys_tmp1081;
	wire signed [31:0] w_sys_tmp1086;
	wire signed [31:0] w_sys_tmp1087;
	wire signed [31:0] w_sys_tmp1092;
	wire signed [31:0] w_sys_tmp1093;
	wire signed [31:0] w_sys_tmp1098;
	wire signed [31:0] w_sys_tmp1099;
	wire signed [31:0] w_sys_tmp1104;
	wire signed [31:0] w_sys_tmp1105;
	wire signed [31:0] w_sys_tmp1110;
	wire signed [31:0] w_sys_tmp1111;
	wire signed [31:0] w_sys_tmp1116;
	wire signed [31:0] w_sys_tmp1117;
	wire signed [31:0] w_sys_tmp1122;
	wire signed [31:0] w_sys_tmp1123;
	wire signed [31:0] w_sys_tmp1128;
	wire signed [31:0] w_sys_tmp1129;
	wire signed [31:0] w_sys_tmp1134;
	wire signed [31:0] w_sys_tmp1135;
	wire signed [31:0] w_sys_tmp1140;
	wire signed [31:0] w_sys_tmp1141;
	wire signed [31:0] w_sys_tmp1146;
	wire signed [31:0] w_sys_tmp1147;
	wire signed [31:0] w_sys_tmp1152;
	wire signed [31:0] w_sys_tmp1153;
	wire signed [31:0] w_sys_tmp1158;
	wire signed [31:0] w_sys_tmp1159;
	wire signed [31:0] w_sys_tmp1164;
	wire signed [31:0] w_sys_tmp1165;
	wire signed [31:0] w_sys_tmp1170;
	wire signed [31:0] w_sys_tmp1171;
	wire signed [31:0] w_sys_tmp1176;
	wire signed [31:0] w_sys_tmp1177;
	wire signed [31:0] w_sys_tmp1182;
	wire signed [31:0] w_sys_tmp1183;
	wire signed [31:0] w_sys_tmp1188;
	wire signed [31:0] w_sys_tmp1189;
	wire signed [31:0] w_sys_tmp1194;
	wire signed [31:0] w_sys_tmp1195;
	wire signed [31:0] w_sys_tmp1200;
	wire signed [31:0] w_sys_tmp1201;
	wire signed [31:0] w_sys_tmp1206;
	wire signed [31:0] w_sys_tmp1207;
	wire signed [31:0] w_sys_tmp1212;
	wire signed [31:0] w_sys_tmp1213;
	wire signed [31:0] w_sys_tmp1218;
	wire signed [31:0] w_sys_tmp1219;
	wire signed [31:0] w_sys_tmp1224;
	wire signed [31:0] w_sys_tmp1225;
	wire signed [31:0] w_sys_tmp1230;
	wire signed [31:0] w_sys_tmp1231;
	wire signed [31:0] w_sys_tmp1236;
	wire signed [31:0] w_sys_tmp1237;
	wire signed [31:0] w_sys_tmp1248;
	wire signed [31:0] w_sys_tmp1249;
	wire signed [31:0] w_sys_tmp1254;
	wire signed [31:0] w_sys_tmp1255;
	wire signed [31:0] w_sys_tmp1266;
	wire signed [31:0] w_sys_tmp1267;
	wire signed [31:0] w_sys_tmp1272;
	wire signed [31:0] w_sys_tmp1273;
	wire signed [31:0] w_sys_tmp1278;
	wire signed [31:0] w_sys_tmp1279;
	wire signed [31:0] w_sys_tmp1284;
	wire signed [31:0] w_sys_tmp1285;
	wire signed [31:0] w_sys_tmp1290;
	wire signed [31:0] w_sys_tmp1291;
	wire signed [31:0] w_sys_tmp1296;
	wire signed [31:0] w_sys_tmp1297;
	wire signed [31:0] w_sys_tmp1302;
	wire signed [31:0] w_sys_tmp1303;
	wire signed [31:0] w_sys_tmp1308;
	wire signed [31:0] w_sys_tmp1309;
	wire signed [31:0] w_sys_tmp1314;
	wire signed [31:0] w_sys_tmp1315;
	wire signed [31:0] w_sys_tmp1320;
	wire signed [31:0] w_sys_tmp1321;
	wire signed [31:0] w_sys_tmp1326;
	wire signed [31:0] w_sys_tmp1327;
	wire signed [31:0] w_sys_tmp1332;
	wire signed [31:0] w_sys_tmp1333;
	wire signed [31:0] w_sys_tmp1338;
	wire signed [31:0] w_sys_tmp1339;
	wire signed [31:0] w_sys_tmp1344;
	wire signed [31:0] w_sys_tmp1345;
	wire signed [31:0] w_sys_tmp1350;
	wire signed [31:0] w_sys_tmp1351;
	wire signed [31:0] w_sys_tmp1356;
	wire signed [31:0] w_sys_tmp1357;
	wire signed [31:0] w_sys_tmp1362;
	wire signed [31:0] w_sys_tmp1363;
	wire signed [31:0] w_sys_tmp1368;
	wire signed [31:0] w_sys_tmp1369;
	wire signed [31:0] w_sys_tmp1374;
	wire signed [31:0] w_sys_tmp1375;
	wire signed [31:0] w_sys_tmp1380;
	wire signed [31:0] w_sys_tmp1381;
	wire signed [31:0] w_sys_tmp1386;
	wire signed [31:0] w_sys_tmp1387;
	wire signed [31:0] w_sys_tmp1392;
	wire signed [31:0] w_sys_tmp1393;
	wire signed [31:0] w_sys_tmp1398;
	wire signed [31:0] w_sys_tmp1399;
	wire signed [31:0] w_sys_tmp1404;
	wire signed [31:0] w_sys_tmp1405;
	wire signed [31:0] w_sys_tmp1410;
	wire signed [31:0] w_sys_tmp1411;
	wire signed [31:0] w_sys_tmp1416;
	wire signed [31:0] w_sys_tmp1417;
	wire signed [31:0] w_sys_tmp1422;
	wire signed [31:0] w_sys_tmp1423;
	wire signed [31:0] w_sys_tmp1428;
	wire signed [31:0] w_sys_tmp1429;
	wire signed [31:0] w_sys_tmp1434;
	wire signed [31:0] w_sys_tmp1435;
	wire signed [31:0] w_sys_tmp1440;
	wire signed [31:0] w_sys_tmp1441;
	wire signed [31:0] w_sys_tmp1446;
	wire signed [31:0] w_sys_tmp1447;
	wire signed [31:0] w_sys_tmp1452;
	wire signed [31:0] w_sys_tmp1453;
	wire signed [31:0] w_sys_tmp1458;
	wire signed [31:0] w_sys_tmp1459;
	wire signed [31:0] w_sys_tmp1464;
	wire signed [31:0] w_sys_tmp1465;
	wire signed [31:0] w_sys_tmp1470;
	wire signed [31:0] w_sys_tmp1471;
	wire signed [31:0] w_sys_tmp1476;
	wire signed [31:0] w_sys_tmp1477;
	wire signed [31:0] w_sys_tmp1482;
	wire signed [31:0] w_sys_tmp1483;
	wire signed [31:0] w_sys_tmp1488;
	wire signed [31:0] w_sys_tmp1489;
	wire signed [31:0] w_sys_tmp1494;
	wire signed [31:0] w_sys_tmp1495;
	wire signed [31:0] w_sys_tmp1500;
	wire signed [31:0] w_sys_tmp1501;
	wire signed [31:0] w_sys_tmp1506;
	wire signed [31:0] w_sys_tmp1507;
	wire signed [31:0] w_sys_tmp1512;
	wire signed [31:0] w_sys_tmp1513;
	wire signed [31:0] w_sys_tmp1518;
	wire signed [31:0] w_sys_tmp1519;
	wire signed [31:0] w_sys_tmp1524;
	wire signed [31:0] w_sys_tmp1525;
	wire signed [31:0] w_sys_tmp1530;
	wire signed [31:0] w_sys_tmp1531;
	wire signed [31:0] w_sys_tmp1536;
	wire signed [31:0] w_sys_tmp1537;
	wire signed [31:0] w_sys_tmp1542;
	wire signed [31:0] w_sys_tmp1543;
	wire signed [31:0] w_sys_tmp1548;
	wire signed [31:0] w_sys_tmp1549;
	wire signed [31:0] w_sys_tmp1554;
	wire signed [31:0] w_sys_tmp1555;
	wire signed [31:0] w_sys_tmp1560;
	wire signed [31:0] w_sys_tmp1561;
	wire signed [31:0] w_sys_tmp1566;
	wire signed [31:0] w_sys_tmp1567;
	wire signed [31:0] w_sys_tmp1572;
	wire signed [31:0] w_sys_tmp1573;
	wire signed [31:0] w_sys_tmp1578;
	wire signed [31:0] w_sys_tmp1579;
	wire signed [31:0] w_sys_tmp1584;
	wire signed [31:0] w_sys_tmp1585;
	wire signed [31:0] w_sys_tmp1590;
	wire signed [31:0] w_sys_tmp1591;
	wire signed [31:0] w_sys_tmp1596;
	wire signed [31:0] w_sys_tmp1597;
	wire signed [31:0] w_sys_tmp1602;
	wire signed [31:0] w_sys_tmp1603;
	wire signed [31:0] w_sys_tmp1608;
	wire signed [31:0] w_sys_tmp1609;
	wire signed [31:0] w_sys_tmp1614;
	wire signed [31:0] w_sys_tmp1615;
	wire signed [31:0] w_sys_tmp1620;
	wire signed [31:0] w_sys_tmp1621;
	wire signed [31:0] w_sys_tmp1626;
	wire signed [31:0] w_sys_tmp1627;
	wire signed [31:0] w_sys_tmp1632;
	wire signed [31:0] w_sys_tmp1633;
	wire signed [31:0] w_sys_tmp1638;
	wire signed [31:0] w_sys_tmp1639;
	wire signed [31:0] w_sys_tmp1644;
	wire signed [31:0] w_sys_tmp1645;
	wire signed [31:0] w_sys_tmp1650;
	wire signed [31:0] w_sys_tmp1651;
	wire signed [31:0] w_sys_tmp1656;
	wire signed [31:0] w_sys_tmp1657;
	wire signed [31:0] w_sys_tmp1662;
	wire signed [31:0] w_sys_tmp1663;
	wire signed [31:0] w_sys_tmp1668;
	wire signed [31:0] w_sys_tmp1669;
	wire signed [31:0] w_sys_tmp1674;
	wire signed [31:0] w_sys_tmp1675;
	wire signed [31:0] w_sys_tmp1680;
	wire signed [31:0] w_sys_tmp1681;
	wire signed [31:0] w_sys_tmp1686;
	wire signed [31:0] w_sys_tmp1687;
	wire signed [31:0] w_sys_tmp1692;
	wire signed [31:0] w_sys_tmp1693;
	wire signed [31:0] w_sys_tmp1698;
	wire signed [31:0] w_sys_tmp1699;
	wire signed [31:0] w_sys_tmp1704;
	wire signed [31:0] w_sys_tmp1705;
	wire signed [31:0] w_sys_tmp1710;
	wire signed [31:0] w_sys_tmp1711;
	wire signed [31:0] w_sys_tmp1716;
	wire signed [31:0] w_sys_tmp1717;
	wire signed [31:0] w_sys_tmp1722;
	wire signed [31:0] w_sys_tmp1723;
	wire signed [31:0] w_sys_tmp1728;
	wire signed [31:0] w_sys_tmp1729;
	wire signed [31:0] w_sys_tmp1734;
	wire signed [31:0] w_sys_tmp1735;
	wire signed [31:0] w_sys_tmp1740;
	wire signed [31:0] w_sys_tmp1741;
	wire signed [31:0] w_sys_tmp1746;
	wire signed [31:0] w_sys_tmp1747;
	wire signed [31:0] w_sys_tmp1752;
	wire signed [31:0] w_sys_tmp1753;
	wire signed [31:0] w_sys_tmp1758;
	wire signed [31:0] w_sys_tmp1759;
	wire signed [31:0] w_sys_tmp1764;
	wire signed [31:0] w_sys_tmp1765;
	wire signed [31:0] w_sys_tmp1770;
	wire signed [31:0] w_sys_tmp1771;
	wire signed [31:0] w_sys_tmp1776;
	wire signed [31:0] w_sys_tmp1777;
	wire signed [31:0] w_sys_tmp1782;
	wire signed [31:0] w_sys_tmp1783;
	wire signed [31:0] w_sys_tmp1788;
	wire signed [31:0] w_sys_tmp1789;
	wire signed [31:0] w_sys_tmp1794;
	wire signed [31:0] w_sys_tmp1795;
	wire signed [31:0] w_sys_tmp1800;
	wire signed [31:0] w_sys_tmp1801;
	wire signed [31:0] w_sys_tmp1806;
	wire signed [31:0] w_sys_tmp1807;
	wire signed [31:0] w_sys_tmp1812;
	wire signed [31:0] w_sys_tmp1813;
	wire signed [31:0] w_sys_tmp1818;
	wire signed [31:0] w_sys_tmp1819;
	wire signed [31:0] w_sys_tmp1824;
	wire signed [31:0] w_sys_tmp1825;
	wire signed [31:0] w_sys_tmp1830;
	wire signed [31:0] w_sys_tmp1831;
	wire signed [31:0] w_sys_tmp1836;
	wire signed [31:0] w_sys_tmp1837;
	wire signed [31:0] w_sys_tmp1842;
	wire signed [31:0] w_sys_tmp1843;
	wire signed [31:0] w_sys_tmp1848;
	wire signed [31:0] w_sys_tmp1849;
	wire signed [31:0] w_sys_tmp1853;
	wire signed [31:0] w_sys_tmp1854;
	wire               w_sys_tmp1855;
	wire               w_sys_tmp1856;
	wire signed [31:0] w_sys_tmp1857;
	wire signed [31:0] w_sys_tmp1860;
	wire signed [31:0] w_sys_tmp1861;
	wire        [31:0] w_sys_tmp1862;
	wire signed [31:0] w_sys_tmp1866;
	wire signed [31:0] w_sys_tmp1867;
	wire signed [31:0] w_sys_tmp1872;
	wire signed [31:0] w_sys_tmp1873;
	wire signed [31:0] w_sys_tmp1878;
	wire signed [31:0] w_sys_tmp1879;
	wire signed [31:0] w_sys_tmp1884;
	wire signed [31:0] w_sys_tmp1885;
	wire signed [31:0] w_sys_tmp1890;
	wire signed [31:0] w_sys_tmp1891;
	wire signed [31:0] w_sys_tmp1896;
	wire signed [31:0] w_sys_tmp1897;
	wire signed [31:0] w_sys_tmp1902;
	wire signed [31:0] w_sys_tmp1903;
	wire signed [31:0] w_sys_tmp1908;
	wire signed [31:0] w_sys_tmp1909;
	wire signed [31:0] w_sys_tmp1914;
	wire signed [31:0] w_sys_tmp1915;
	wire signed [31:0] w_sys_tmp1920;
	wire signed [31:0] w_sys_tmp1921;
	wire signed [31:0] w_sys_tmp1926;
	wire signed [31:0] w_sys_tmp1927;
	wire signed [31:0] w_sys_tmp1932;
	wire signed [31:0] w_sys_tmp1933;
	wire signed [31:0] w_sys_tmp1938;
	wire signed [31:0] w_sys_tmp1939;
	wire signed [31:0] w_sys_tmp1944;
	wire signed [31:0] w_sys_tmp1945;
	wire signed [31:0] w_sys_tmp1950;
	wire signed [31:0] w_sys_tmp1951;
	wire signed [31:0] w_sys_tmp1956;
	wire signed [31:0] w_sys_tmp1957;
	wire signed [31:0] w_sys_tmp1962;
	wire signed [31:0] w_sys_tmp1963;
	wire signed [31:0] w_sys_tmp1968;
	wire signed [31:0] w_sys_tmp1969;
	wire signed [31:0] w_sys_tmp1974;
	wire signed [31:0] w_sys_tmp1975;
	wire signed [31:0] w_sys_tmp1980;
	wire signed [31:0] w_sys_tmp1981;
	wire signed [31:0] w_sys_tmp1986;
	wire signed [31:0] w_sys_tmp1987;
	wire signed [31:0] w_sys_tmp1992;
	wire signed [31:0] w_sys_tmp1993;
	wire signed [31:0] w_sys_tmp1998;
	wire signed [31:0] w_sys_tmp1999;
	wire signed [31:0] w_sys_tmp2004;
	wire signed [31:0] w_sys_tmp2005;
	wire signed [31:0] w_sys_tmp2010;
	wire signed [31:0] w_sys_tmp2011;
	wire signed [31:0] w_sys_tmp2016;
	wire signed [31:0] w_sys_tmp2017;
	wire signed [31:0] w_sys_tmp2022;
	wire signed [31:0] w_sys_tmp2023;
	wire signed [31:0] w_sys_tmp2028;
	wire signed [31:0] w_sys_tmp2029;
	wire signed [31:0] w_sys_tmp2034;
	wire signed [31:0] w_sys_tmp2035;
	wire signed [31:0] w_sys_tmp2040;
	wire signed [31:0] w_sys_tmp2041;
	wire signed [31:0] w_sys_tmp2046;
	wire signed [31:0] w_sys_tmp2047;
	wire signed [31:0] w_sys_tmp2051;
	wire signed [31:0] w_sys_tmp2052;
	wire signed [31:0] w_sys_tmp2056;
	wire signed [31:0] w_sys_tmp2057;
	wire signed [31:0] w_sys_tmp2061;
	wire signed [31:0] w_sys_tmp2062;
	wire signed [31:0] w_sys_tmp2066;
	wire signed [31:0] w_sys_tmp2067;
	wire signed [31:0] w_sys_tmp2071;
	wire signed [31:0] w_sys_tmp2072;
	wire signed [31:0] w_sys_tmp2076;
	wire signed [31:0] w_sys_tmp2077;
	wire signed [31:0] w_sys_tmp2081;
	wire signed [31:0] w_sys_tmp2082;
	wire signed [31:0] w_sys_tmp2086;
	wire signed [31:0] w_sys_tmp2087;
	wire signed [31:0] w_sys_tmp2091;
	wire signed [31:0] w_sys_tmp2092;
	wire signed [31:0] w_sys_tmp2096;
	wire signed [31:0] w_sys_tmp2097;
	wire signed [31:0] w_sys_tmp2101;
	wire signed [31:0] w_sys_tmp2102;
	wire signed [31:0] w_sys_tmp2106;
	wire signed [31:0] w_sys_tmp2107;
	wire signed [31:0] w_sys_tmp2111;
	wire signed [31:0] w_sys_tmp2112;
	wire signed [31:0] w_sys_tmp2116;
	wire signed [31:0] w_sys_tmp2117;
	wire signed [31:0] w_sys_tmp2121;
	wire signed [31:0] w_sys_tmp2122;
	wire signed [31:0] w_sys_tmp2126;
	wire signed [31:0] w_sys_tmp2127;
	wire signed [31:0] w_sys_tmp2131;
	wire signed [31:0] w_sys_tmp2132;
	wire signed [31:0] w_sys_tmp2136;
	wire signed [31:0] w_sys_tmp2137;
	wire signed [31:0] w_sys_tmp2141;
	wire signed [31:0] w_sys_tmp2142;
	wire signed [31:0] w_sys_tmp2146;
	wire signed [31:0] w_sys_tmp2147;
	wire signed [31:0] w_sys_tmp2151;
	wire signed [31:0] w_sys_tmp2152;
	wire signed [31:0] w_sys_tmp2156;
	wire signed [31:0] w_sys_tmp2157;
	wire signed [31:0] w_sys_tmp2161;
	wire signed [31:0] w_sys_tmp2162;
	wire signed [31:0] w_sys_tmp2166;
	wire signed [31:0] w_sys_tmp2167;
	wire signed [31:0] w_sys_tmp2171;
	wire signed [31:0] w_sys_tmp2172;
	wire signed [31:0] w_sys_tmp2176;
	wire signed [31:0] w_sys_tmp2177;
	wire signed [31:0] w_sys_tmp2181;
	wire signed [31:0] w_sys_tmp2182;
	wire signed [31:0] w_sys_tmp2186;
	wire signed [31:0] w_sys_tmp2187;
	wire signed [31:0] w_sys_tmp2191;
	wire signed [31:0] w_sys_tmp2192;
	wire signed [31:0] w_sys_tmp2196;
	wire signed [31:0] w_sys_tmp2197;
	wire signed [31:0] w_sys_tmp2201;
	wire signed [31:0] w_sys_tmp2202;
	wire signed [31:0] w_sys_tmp2206;
	wire signed [31:0] w_sys_tmp2207;
	wire signed [31:0] w_sys_tmp2211;
	wire signed [31:0] w_sys_tmp2212;
	wire signed [31:0] w_sys_tmp2216;
	wire signed [31:0] w_sys_tmp2217;
	wire signed [31:0] w_sys_tmp2221;
	wire signed [31:0] w_sys_tmp2222;
	wire signed [31:0] w_sys_tmp2226;
	wire signed [31:0] w_sys_tmp2227;
	wire signed [31:0] w_sys_tmp2231;
	wire signed [31:0] w_sys_tmp2232;
	wire signed [31:0] w_sys_tmp2236;
	wire signed [31:0] w_sys_tmp2237;
	wire signed [31:0] w_sys_tmp2241;
	wire signed [31:0] w_sys_tmp2242;
	wire signed [31:0] w_sys_tmp2246;
	wire signed [31:0] w_sys_tmp2247;
	wire signed [31:0] w_sys_tmp2251;
	wire signed [31:0] w_sys_tmp2252;
	wire signed [31:0] w_sys_tmp2256;
	wire signed [31:0] w_sys_tmp2257;
	wire signed [31:0] w_sys_tmp2261;
	wire signed [31:0] w_sys_tmp2262;
	wire signed [31:0] w_sys_tmp2266;
	wire signed [31:0] w_sys_tmp2267;
	wire signed [31:0] w_sys_tmp2271;
	wire signed [31:0] w_sys_tmp2272;
	wire signed [31:0] w_sys_tmp2276;
	wire signed [31:0] w_sys_tmp2277;
	wire signed [31:0] w_sys_tmp2281;
	wire signed [31:0] w_sys_tmp2282;
	wire signed [31:0] w_sys_tmp2286;
	wire signed [31:0] w_sys_tmp2287;
	wire signed [31:0] w_sys_tmp2291;
	wire signed [31:0] w_sys_tmp2292;
	wire signed [31:0] w_sys_tmp2296;
	wire signed [31:0] w_sys_tmp2297;
	wire signed [31:0] w_sys_tmp2301;
	wire signed [31:0] w_sys_tmp2302;
	wire signed [31:0] w_sys_tmp2306;
	wire signed [31:0] w_sys_tmp2307;
	wire signed [31:0] w_sys_tmp2311;
	wire signed [31:0] w_sys_tmp2312;
	wire signed [31:0] w_sys_tmp2316;
	wire signed [31:0] w_sys_tmp2317;
	wire signed [31:0] w_sys_tmp2321;
	wire signed [31:0] w_sys_tmp2322;
	wire signed [31:0] w_sys_tmp2326;
	wire signed [31:0] w_sys_tmp2327;
	wire signed [31:0] w_sys_tmp2331;
	wire signed [31:0] w_sys_tmp2332;
	wire signed [31:0] w_sys_tmp2336;
	wire signed [31:0] w_sys_tmp2337;
	wire signed [31:0] w_sys_tmp2341;
	wire signed [31:0] w_sys_tmp2342;
	wire signed [31:0] w_sys_tmp2346;
	wire signed [31:0] w_sys_tmp2347;
	wire signed [31:0] w_sys_tmp2351;
	wire signed [31:0] w_sys_tmp2352;
	wire signed [31:0] w_sys_tmp2356;
	wire signed [31:0] w_sys_tmp2357;
	wire signed [31:0] w_sys_tmp2361;
	wire signed [31:0] w_sys_tmp2362;
	wire signed [31:0] w_sys_tmp2366;
	wire signed [31:0] w_sys_tmp2367;
	wire signed [31:0] w_sys_tmp2371;
	wire signed [31:0] w_sys_tmp2372;
	wire signed [31:0] w_sys_tmp2376;
	wire signed [31:0] w_sys_tmp2377;
	wire signed [31:0] w_sys_tmp2381;
	wire signed [31:0] w_sys_tmp2382;
	wire signed [31:0] w_sys_tmp2386;
	wire signed [31:0] w_sys_tmp2387;
	wire signed [31:0] w_sys_tmp2391;
	wire signed [31:0] w_sys_tmp2392;
	wire signed [31:0] w_sys_tmp2396;
	wire signed [31:0] w_sys_tmp2397;
	wire signed [31:0] w_sys_tmp2401;
	wire signed [31:0] w_sys_tmp2402;
	wire signed [31:0] w_sys_tmp2406;
	wire signed [31:0] w_sys_tmp2407;
	wire signed [31:0] w_sys_tmp2411;
	wire signed [31:0] w_sys_tmp2412;
	wire signed [31:0] w_sys_tmp2416;
	wire signed [31:0] w_sys_tmp2417;
	wire signed [31:0] w_sys_tmp2421;
	wire signed [31:0] w_sys_tmp2422;
	wire signed [31:0] w_sys_tmp2426;
	wire signed [31:0] w_sys_tmp2427;
	wire signed [31:0] w_sys_tmp2431;
	wire signed [31:0] w_sys_tmp2432;
	wire signed [31:0] w_sys_tmp2436;
	wire signed [31:0] w_sys_tmp2437;
	wire signed [31:0] w_sys_tmp2441;
	wire signed [31:0] w_sys_tmp2442;
	wire signed [31:0] w_sys_tmp2446;
	wire signed [31:0] w_sys_tmp2447;
	wire signed [31:0] w_sys_tmp2451;
	wire signed [31:0] w_sys_tmp2452;
	wire signed [31:0] w_sys_tmp2456;
	wire signed [31:0] w_sys_tmp2457;
	wire signed [31:0] w_sys_tmp2461;
	wire signed [31:0] w_sys_tmp2462;
	wire signed [31:0] w_sys_tmp2466;
	wire signed [31:0] w_sys_tmp2467;
	wire signed [31:0] w_sys_tmp2471;
	wire signed [31:0] w_sys_tmp2472;
	wire signed [31:0] w_sys_tmp2476;
	wire signed [31:0] w_sys_tmp2477;
	wire signed [31:0] w_sys_tmp2481;
	wire signed [31:0] w_sys_tmp2482;
	wire signed [31:0] w_sys_tmp2486;
	wire signed [31:0] w_sys_tmp2487;
	wire signed [31:0] w_sys_tmp2491;
	wire signed [31:0] w_sys_tmp2492;
	wire signed [31:0] w_sys_tmp2496;
	wire signed [31:0] w_sys_tmp2497;
	wire signed [31:0] w_sys_tmp2501;
	wire signed [31:0] w_sys_tmp2502;
	wire signed [31:0] w_sys_tmp2506;
	wire signed [31:0] w_sys_tmp2507;
	wire signed [31:0] w_sys_tmp2511;
	wire signed [31:0] w_sys_tmp2512;
	wire signed [31:0] w_sys_tmp2516;
	wire signed [31:0] w_sys_tmp2517;
	wire signed [31:0] w_sys_tmp2521;
	wire signed [31:0] w_sys_tmp2522;
	wire signed [31:0] w_sys_tmp2525;
	wire signed [31:0] w_sys_tmp2526;
	wire               w_sys_tmp2527;
	wire               w_sys_tmp2528;
	wire signed [31:0] w_sys_tmp2529;
	wire signed [31:0] w_sys_tmp2532;
	wire signed [31:0] w_sys_tmp2533;
	wire        [31:0] w_sys_tmp2534;
	wire signed [31:0] w_sys_tmp2538;
	wire signed [31:0] w_sys_tmp2539;
	wire signed [31:0] w_sys_tmp2544;
	wire signed [31:0] w_sys_tmp2545;
	wire signed [31:0] w_sys_tmp2550;
	wire signed [31:0] w_sys_tmp2551;
	wire signed [31:0] w_sys_tmp2556;
	wire signed [31:0] w_sys_tmp2557;
	wire signed [31:0] w_sys_tmp2562;
	wire signed [31:0] w_sys_tmp2563;
	wire signed [31:0] w_sys_tmp2568;
	wire signed [31:0] w_sys_tmp2569;
	wire signed [31:0] w_sys_tmp2574;
	wire signed [31:0] w_sys_tmp2575;
	wire signed [31:0] w_sys_tmp2580;
	wire signed [31:0] w_sys_tmp2581;
	wire signed [31:0] w_sys_tmp2586;
	wire signed [31:0] w_sys_tmp2587;
	wire signed [31:0] w_sys_tmp2592;
	wire signed [31:0] w_sys_tmp2593;
	wire signed [31:0] w_sys_tmp2598;
	wire signed [31:0] w_sys_tmp2599;
	wire signed [31:0] w_sys_tmp2604;
	wire signed [31:0] w_sys_tmp2605;
	wire signed [31:0] w_sys_tmp2610;
	wire signed [31:0] w_sys_tmp2611;
	wire signed [31:0] w_sys_tmp2616;
	wire signed [31:0] w_sys_tmp2617;
	wire signed [31:0] w_sys_tmp2622;
	wire signed [31:0] w_sys_tmp2623;
	wire signed [31:0] w_sys_tmp2628;
	wire signed [31:0] w_sys_tmp2629;
	wire signed [31:0] w_sys_tmp2634;
	wire signed [31:0] w_sys_tmp2635;
	wire signed [31:0] w_sys_tmp2640;
	wire signed [31:0] w_sys_tmp2641;
	wire signed [31:0] w_sys_tmp2646;
	wire signed [31:0] w_sys_tmp2647;
	wire signed [31:0] w_sys_tmp2652;
	wire signed [31:0] w_sys_tmp2653;
	wire signed [31:0] w_sys_tmp2658;
	wire signed [31:0] w_sys_tmp2659;
	wire signed [31:0] w_sys_tmp2664;
	wire signed [31:0] w_sys_tmp2665;
	wire signed [31:0] w_sys_tmp2670;
	wire signed [31:0] w_sys_tmp2671;
	wire signed [31:0] w_sys_tmp2676;
	wire signed [31:0] w_sys_tmp2677;
	wire signed [31:0] w_sys_tmp2682;
	wire signed [31:0] w_sys_tmp2683;
	wire signed [31:0] w_sys_tmp2688;
	wire signed [31:0] w_sys_tmp2689;
	wire signed [31:0] w_sys_tmp2694;
	wire signed [31:0] w_sys_tmp2695;
	wire signed [31:0] w_sys_tmp2700;
	wire signed [31:0] w_sys_tmp2701;
	wire signed [31:0] w_sys_tmp2706;
	wire signed [31:0] w_sys_tmp2707;
	wire signed [31:0] w_sys_tmp2712;
	wire signed [31:0] w_sys_tmp2713;
	wire signed [31:0] w_sys_tmp2718;
	wire signed [31:0] w_sys_tmp2719;
	wire signed [31:0] w_sys_tmp2723;
	wire signed [31:0] w_sys_tmp2724;
	wire signed [31:0] w_sys_tmp2728;
	wire signed [31:0] w_sys_tmp2729;
	wire signed [31:0] w_sys_tmp2733;
	wire signed [31:0] w_sys_tmp2734;
	wire signed [31:0] w_sys_tmp2738;
	wire signed [31:0] w_sys_tmp2739;
	wire signed [31:0] w_sys_tmp2743;
	wire signed [31:0] w_sys_tmp2744;
	wire signed [31:0] w_sys_tmp2748;
	wire signed [31:0] w_sys_tmp2749;
	wire signed [31:0] w_sys_tmp2753;
	wire signed [31:0] w_sys_tmp2754;
	wire signed [31:0] w_sys_tmp2758;
	wire signed [31:0] w_sys_tmp2759;
	wire signed [31:0] w_sys_tmp2763;
	wire signed [31:0] w_sys_tmp2764;
	wire signed [31:0] w_sys_tmp2768;
	wire signed [31:0] w_sys_tmp2769;
	wire signed [31:0] w_sys_tmp2773;
	wire signed [31:0] w_sys_tmp2774;
	wire signed [31:0] w_sys_tmp2778;
	wire signed [31:0] w_sys_tmp2779;
	wire signed [31:0] w_sys_tmp2783;
	wire signed [31:0] w_sys_tmp2784;
	wire signed [31:0] w_sys_tmp2788;
	wire signed [31:0] w_sys_tmp2789;
	wire signed [31:0] w_sys_tmp2793;
	wire signed [31:0] w_sys_tmp2794;
	wire signed [31:0] w_sys_tmp2798;
	wire signed [31:0] w_sys_tmp2799;
	wire signed [31:0] w_sys_tmp2803;
	wire signed [31:0] w_sys_tmp2804;
	wire signed [31:0] w_sys_tmp2808;
	wire signed [31:0] w_sys_tmp2809;
	wire signed [31:0] w_sys_tmp2813;
	wire signed [31:0] w_sys_tmp2814;
	wire signed [31:0] w_sys_tmp2818;
	wire signed [31:0] w_sys_tmp2819;
	wire signed [31:0] w_sys_tmp2823;
	wire signed [31:0] w_sys_tmp2824;
	wire signed [31:0] w_sys_tmp2828;
	wire signed [31:0] w_sys_tmp2829;
	wire signed [31:0] w_sys_tmp2833;
	wire signed [31:0] w_sys_tmp2834;
	wire signed [31:0] w_sys_tmp2838;
	wire signed [31:0] w_sys_tmp2839;
	wire signed [31:0] w_sys_tmp2843;
	wire signed [31:0] w_sys_tmp2844;
	wire signed [31:0] w_sys_tmp2848;
	wire signed [31:0] w_sys_tmp2849;
	wire signed [31:0] w_sys_tmp2853;
	wire signed [31:0] w_sys_tmp2854;
	wire signed [31:0] w_sys_tmp2858;
	wire signed [31:0] w_sys_tmp2859;
	wire signed [31:0] w_sys_tmp2863;
	wire signed [31:0] w_sys_tmp2864;
	wire signed [31:0] w_sys_tmp2868;
	wire signed [31:0] w_sys_tmp2869;
	wire signed [31:0] w_sys_tmp2873;
	wire signed [31:0] w_sys_tmp2874;
	wire signed [31:0] w_sys_tmp2878;
	wire signed [31:0] w_sys_tmp2879;
	wire signed [31:0] w_sys_tmp2883;
	wire signed [31:0] w_sys_tmp2884;
	wire signed [31:0] w_sys_tmp2888;
	wire signed [31:0] w_sys_tmp2889;
	wire signed [31:0] w_sys_tmp2893;
	wire signed [31:0] w_sys_tmp2894;
	wire signed [31:0] w_sys_tmp2898;
	wire signed [31:0] w_sys_tmp2899;
	wire signed [31:0] w_sys_tmp2903;
	wire signed [31:0] w_sys_tmp2904;
	wire signed [31:0] w_sys_tmp2908;
	wire signed [31:0] w_sys_tmp2909;
	wire signed [31:0] w_sys_tmp2913;
	wire signed [31:0] w_sys_tmp2914;
	wire signed [31:0] w_sys_tmp2918;
	wire signed [31:0] w_sys_tmp2919;
	wire signed [31:0] w_sys_tmp2923;
	wire signed [31:0] w_sys_tmp2924;
	wire signed [31:0] w_sys_tmp2928;
	wire signed [31:0] w_sys_tmp2929;
	wire signed [31:0] w_sys_tmp2933;
	wire signed [31:0] w_sys_tmp2934;
	wire signed [31:0] w_sys_tmp2938;
	wire signed [31:0] w_sys_tmp2939;
	wire signed [31:0] w_sys_tmp2943;
	wire signed [31:0] w_sys_tmp2944;
	wire signed [31:0] w_sys_tmp2948;
	wire signed [31:0] w_sys_tmp2949;
	wire signed [31:0] w_sys_tmp2953;
	wire signed [31:0] w_sys_tmp2954;
	wire signed [31:0] w_sys_tmp2958;
	wire signed [31:0] w_sys_tmp2959;
	wire signed [31:0] w_sys_tmp2963;
	wire signed [31:0] w_sys_tmp2964;
	wire signed [31:0] w_sys_tmp2968;
	wire signed [31:0] w_sys_tmp2969;
	wire signed [31:0] w_sys_tmp2973;
	wire signed [31:0] w_sys_tmp2974;
	wire signed [31:0] w_sys_tmp2978;
	wire signed [31:0] w_sys_tmp2979;
	wire signed [31:0] w_sys_tmp2983;
	wire signed [31:0] w_sys_tmp2984;
	wire signed [31:0] w_sys_tmp2988;
	wire signed [31:0] w_sys_tmp2989;
	wire signed [31:0] w_sys_tmp2993;
	wire signed [31:0] w_sys_tmp2994;
	wire signed [31:0] w_sys_tmp2998;
	wire signed [31:0] w_sys_tmp2999;
	wire signed [31:0] w_sys_tmp3003;
	wire signed [31:0] w_sys_tmp3004;
	wire signed [31:0] w_sys_tmp3008;
	wire signed [31:0] w_sys_tmp3009;
	wire signed [31:0] w_sys_tmp3013;
	wire signed [31:0] w_sys_tmp3014;
	wire signed [31:0] w_sys_tmp3018;
	wire signed [31:0] w_sys_tmp3019;
	wire signed [31:0] w_sys_tmp3023;
	wire signed [31:0] w_sys_tmp3024;
	wire signed [31:0] w_sys_tmp3028;
	wire signed [31:0] w_sys_tmp3029;
	wire signed [31:0] w_sys_tmp3033;
	wire signed [31:0] w_sys_tmp3034;
	wire signed [31:0] w_sys_tmp3038;
	wire signed [31:0] w_sys_tmp3039;
	wire signed [31:0] w_sys_tmp3043;
	wire signed [31:0] w_sys_tmp3044;
	wire signed [31:0] w_sys_tmp3048;
	wire signed [31:0] w_sys_tmp3049;
	wire signed [31:0] w_sys_tmp3053;
	wire signed [31:0] w_sys_tmp3054;
	wire signed [31:0] w_sys_tmp3058;
	wire signed [31:0] w_sys_tmp3059;
	wire signed [31:0] w_sys_tmp3063;
	wire signed [31:0] w_sys_tmp3064;
	wire signed [31:0] w_sys_tmp3068;
	wire signed [31:0] w_sys_tmp3069;
	wire signed [31:0] w_sys_tmp3073;
	wire signed [31:0] w_sys_tmp3074;
	wire signed [31:0] w_sys_tmp3078;
	wire signed [31:0] w_sys_tmp3079;
	wire signed [31:0] w_sys_tmp3083;
	wire signed [31:0] w_sys_tmp3084;
	wire signed [31:0] w_sys_tmp3088;
	wire signed [31:0] w_sys_tmp3089;
	wire signed [31:0] w_sys_tmp3093;
	wire signed [31:0] w_sys_tmp3094;
	wire signed [31:0] w_sys_tmp3098;
	wire signed [31:0] w_sys_tmp3099;
	wire signed [31:0] w_sys_tmp3103;
	wire signed [31:0] w_sys_tmp3104;
	wire signed [31:0] w_sys_tmp3108;
	wire signed [31:0] w_sys_tmp3109;
	wire signed [31:0] w_sys_tmp3113;
	wire signed [31:0] w_sys_tmp3114;
	wire signed [31:0] w_sys_tmp3118;
	wire signed [31:0] w_sys_tmp3119;
	wire signed [31:0] w_sys_tmp3123;
	wire signed [31:0] w_sys_tmp3124;
	wire signed [31:0] w_sys_tmp3128;
	wire signed [31:0] w_sys_tmp3129;
	wire signed [31:0] w_sys_tmp3133;
	wire signed [31:0] w_sys_tmp3134;
	wire signed [31:0] w_sys_tmp3138;
	wire signed [31:0] w_sys_tmp3139;
	wire signed [31:0] w_sys_tmp3143;
	wire signed [31:0] w_sys_tmp3144;
	wire signed [31:0] w_sys_tmp3148;
	wire signed [31:0] w_sys_tmp3149;
	wire signed [31:0] w_sys_tmp3153;
	wire signed [31:0] w_sys_tmp3154;
	wire signed [31:0] w_sys_tmp3158;
	wire signed [31:0] w_sys_tmp3159;
	wire signed [31:0] w_sys_tmp3163;
	wire signed [31:0] w_sys_tmp3164;
	wire signed [31:0] w_sys_tmp3168;
	wire signed [31:0] w_sys_tmp3169;
	wire signed [31:0] w_sys_tmp3173;
	wire signed [31:0] w_sys_tmp3174;
	wire signed [31:0] w_sys_tmp3178;
	wire signed [31:0] w_sys_tmp3179;
	wire signed [31:0] w_sys_tmp3183;
	wire signed [31:0] w_sys_tmp3184;
	wire signed [31:0] w_sys_tmp3188;
	wire signed [31:0] w_sys_tmp3189;
	wire signed [31:0] w_sys_tmp3193;
	wire signed [31:0] w_sys_tmp3194;
	wire signed [31:0] w_sys_tmp3197;
	wire        [31:0] w_sys_tmp3198;
	wire signed [31:0] w_sys_tmp3199;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign o_run_return = r_sys_run_return;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 4'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 8'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 15'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 15'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 15'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 15'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 15'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 15'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 15'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 15'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 15'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 15'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 15'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 15'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 15'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 15'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 15'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 15'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = 32'h3c000000;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'h4103126f;
	assign w_sys_tmp8 = ( !w_sys_tmp9 );
	assign w_sys_tmp9 = (r_run_my_13 < r_run_k_9);
	assign w_sys_tmp10 = (r_run_k_9 + w_sys_intOne);
	assign w_sys_tmp11 = ( !w_sys_tmp12 );
	assign w_sys_tmp12 = (r_run_mx_12 < r_run_j_10);
	assign w_sys_tmp15 = (w_sys_tmp16 + r_run_k_9);
	assign w_sys_tmp16 = (r_run_j_10 * w_sys_tmp17);
	assign w_sys_tmp17 = 32'sh00000081;
	assign w_sys_tmp18 = 32'h0;
	assign w_sys_tmp19 = (r_run_j_10 + w_sys_intOne);
	assign w_sys_tmp56 = ( !w_sys_tmp57 );
	assign w_sys_tmp57 = (r_run_nlast_14 < r_run_n_11);
	assign w_sys_tmp58 = (r_run_n_11 + w_sys_intOne);
	assign w_sys_tmp59 = ( !w_sys_tmp60 );
	assign w_sys_tmp60 = (r_run_my_13 < r_run_j_10);
	assign w_sys_tmp63 = (w_sys_tmp64 + r_run_j_10);
	assign w_sys_tmp64 = 32'sh00000081;
	assign w_sys_tmp65 = 32'h3f000000;
	assign w_sys_tmp67 = (w_sys_tmp68 + r_run_copy2_j_22);
	assign w_sys_tmp68 = (r_run_mx_12 * w_sys_tmp64);
	assign w_sys_tmp70 = 32'h0;
	assign w_sys_tmp72 = (w_sys_tmp73 + w_sys_intOne);
	assign w_sys_tmp73 = (r_run_copy1_j_21 * w_sys_tmp64);
	assign w_sys_tmp75 = 32'h3f800000;
	assign w_sys_tmp77 = (w_sys_tmp78 + r_run_my_13);
	assign w_sys_tmp78 = (r_run_copy0_j_20 * w_sys_tmp79);
	assign w_sys_tmp79 = 32'sh00000015;
	assign w_sys_tmp81 = (r_run_copy0_j_20 + w_sys_intOne);
	assign w_sys_tmp82 = (r_run_copy1_j_21 + w_sys_intOne);
	assign w_sys_tmp83 = (r_run_copy2_j_22 + w_sys_intOne);
	assign w_sys_tmp84 = (r_run_j_10 + w_sys_intOne);
	assign w_sys_tmp223 = ( !w_sys_tmp224 );
	assign w_sys_tmp224 = (w_sys_tmp225 < r_run_k_9);
	assign w_sys_tmp225 = 32'sh00000041;
	assign w_sys_tmp228 = (w_sys_tmp229 + r_run_k_9);
	assign w_sys_tmp229 = 32'sh00000081;
	assign w_sys_tmp230 = w_fld_u_0_dataout_1;
	assign w_sys_tmp234 = (w_sys_tmp235 + r_run_k_9);
	assign w_sys_tmp235 = 32'sh00000102;
	assign w_sys_tmp240 = (w_sys_tmp241 + r_run_k_9);
	assign w_sys_tmp241 = 32'sh00000183;
	assign w_sys_tmp246 = (w_sys_tmp247 + r_run_k_9);
	assign w_sys_tmp247 = 32'sh00000204;
	assign w_sys_tmp252 = (w_sys_tmp253 + r_run_k_9);
	assign w_sys_tmp253 = 32'sh00000285;
	assign w_sys_tmp258 = (w_sys_tmp259 + r_run_k_9);
	assign w_sys_tmp259 = 32'sh00000306;
	assign w_sys_tmp264 = (w_sys_tmp265 + r_run_k_9);
	assign w_sys_tmp265 = 32'sh00000387;
	assign w_sys_tmp270 = (w_sys_tmp271 + r_run_k_9);
	assign w_sys_tmp271 = 32'sh00000408;
	assign w_sys_tmp276 = (w_sys_tmp277 + r_run_k_9);
	assign w_sys_tmp277 = 32'sh00000489;
	assign w_sys_tmp282 = (w_sys_tmp283 + r_run_k_9);
	assign w_sys_tmp283 = 32'sh0000050a;
	assign w_sys_tmp288 = (w_sys_tmp289 + r_run_k_9);
	assign w_sys_tmp289 = 32'sh0000058b;
	assign w_sys_tmp294 = (w_sys_tmp295 + r_run_k_9);
	assign w_sys_tmp295 = 32'sh0000060c;
	assign w_sys_tmp300 = (w_sys_tmp301 + r_run_k_9);
	assign w_sys_tmp301 = 32'sh0000068d;
	assign w_sys_tmp306 = (w_sys_tmp307 + r_run_k_9);
	assign w_sys_tmp307 = 32'sh0000070e;
	assign w_sys_tmp312 = (w_sys_tmp313 + r_run_k_9);
	assign w_sys_tmp313 = 32'sh0000078f;
	assign w_sys_tmp318 = (w_sys_tmp319 + r_run_k_9);
	assign w_sys_tmp319 = 32'sh00000810;
	assign w_sys_tmp324 = (w_sys_tmp325 + r_run_k_9);
	assign w_sys_tmp325 = 32'sh00000891;
	assign w_sys_tmp330 = (w_sys_tmp331 + r_run_k_9);
	assign w_sys_tmp331 = 32'sh00000912;
	assign w_sys_tmp336 = (w_sys_tmp337 + r_run_k_9);
	assign w_sys_tmp337 = 32'sh00000993;
	assign w_sys_tmp342 = (w_sys_tmp343 + r_run_k_9);
	assign w_sys_tmp343 = 32'sh00000a14;
	assign w_sys_tmp348 = (w_sys_tmp349 + r_run_k_9);
	assign w_sys_tmp349 = 32'sh00000a95;
	assign w_sys_tmp354 = (w_sys_tmp355 + r_run_k_9);
	assign w_sys_tmp355 = 32'sh00000b16;
	assign w_sys_tmp360 = (w_sys_tmp361 + r_run_k_9);
	assign w_sys_tmp361 = 32'sh00000b97;
	assign w_sys_tmp366 = (w_sys_tmp367 + r_run_k_9);
	assign w_sys_tmp367 = 32'sh00000c18;
	assign w_sys_tmp372 = (w_sys_tmp373 + r_run_k_9);
	assign w_sys_tmp373 = 32'sh00000c99;
	assign w_sys_tmp378 = (w_sys_tmp379 + r_run_k_9);
	assign w_sys_tmp379 = 32'sh00000d1a;
	assign w_sys_tmp384 = (w_sys_tmp385 + r_run_k_9);
	assign w_sys_tmp385 = 32'sh00000d9b;
	assign w_sys_tmp390 = (w_sys_tmp391 + r_run_k_9);
	assign w_sys_tmp391 = 32'sh00000e1c;
	assign w_sys_tmp396 = (w_sys_tmp397 + r_run_k_9);
	assign w_sys_tmp397 = 32'sh00000e9d;
	assign w_sys_tmp402 = (w_sys_tmp403 + r_run_k_9);
	assign w_sys_tmp403 = 32'sh00000f1e;
	assign w_sys_tmp408 = (w_sys_tmp409 + r_run_k_9);
	assign w_sys_tmp409 = 32'sh00000f9f;
	assign w_sys_tmp414 = (w_sys_tmp415 + r_run_k_9);
	assign w_sys_tmp415 = 32'sh00001020;
	assign w_sys_tmp420 = (w_sys_tmp421 + r_run_k_9);
	assign w_sys_tmp421 = 32'sh000010a1;
	assign w_sys_tmp432 = (w_sys_tmp433 + r_run_k_9);
	assign w_sys_tmp433 = 32'sh00001040;
	assign w_sys_tmp438 = (w_sys_tmp439 + r_run_k_9);
	assign w_sys_tmp439 = 32'sh00001060;
	assign w_sys_tmp450 = (w_sys_tmp451 + r_run_k_9);
	assign w_sys_tmp451 = 32'sh000010c1;
	assign w_sys_tmp456 = (w_sys_tmp457 + r_run_k_9);
	assign w_sys_tmp457 = 32'sh000010e1;
	assign w_sys_tmp462 = (w_sys_tmp463 + r_run_k_9);
	assign w_sys_tmp463 = 32'sh00001122;
	assign w_sys_tmp468 = (w_sys_tmp469 + r_run_k_9);
	assign w_sys_tmp469 = 32'sh00001142;
	assign w_sys_tmp474 = (w_sys_tmp475 + r_run_k_9);
	assign w_sys_tmp475 = 32'sh00001162;
	assign w_sys_tmp480 = (w_sys_tmp481 + r_run_k_9);
	assign w_sys_tmp481 = 32'sh000011a3;
	assign w_sys_tmp486 = (w_sys_tmp487 + r_run_k_9);
	assign w_sys_tmp487 = 32'sh000011c3;
	assign w_sys_tmp492 = (w_sys_tmp493 + r_run_k_9);
	assign w_sys_tmp493 = 32'sh000011e3;
	assign w_sys_tmp498 = (w_sys_tmp499 + r_run_k_9);
	assign w_sys_tmp499 = 32'sh00001224;
	assign w_sys_tmp504 = (w_sys_tmp505 + r_run_k_9);
	assign w_sys_tmp505 = 32'sh00001244;
	assign w_sys_tmp510 = (w_sys_tmp511 + r_run_k_9);
	assign w_sys_tmp511 = 32'sh00001264;
	assign w_sys_tmp516 = (w_sys_tmp517 + r_run_k_9);
	assign w_sys_tmp517 = 32'sh000012a5;
	assign w_sys_tmp522 = (w_sys_tmp523 + r_run_k_9);
	assign w_sys_tmp523 = 32'sh000012c5;
	assign w_sys_tmp528 = (w_sys_tmp529 + r_run_k_9);
	assign w_sys_tmp529 = 32'sh000012e5;
	assign w_sys_tmp534 = (w_sys_tmp535 + r_run_k_9);
	assign w_sys_tmp535 = 32'sh00001326;
	assign w_sys_tmp540 = (w_sys_tmp541 + r_run_k_9);
	assign w_sys_tmp541 = 32'sh00001346;
	assign w_sys_tmp546 = (w_sys_tmp547 + r_run_k_9);
	assign w_sys_tmp547 = 32'sh00001366;
	assign w_sys_tmp552 = (w_sys_tmp553 + r_run_k_9);
	assign w_sys_tmp553 = 32'sh000013a7;
	assign w_sys_tmp558 = (w_sys_tmp559 + r_run_k_9);
	assign w_sys_tmp559 = 32'sh000013c7;
	assign w_sys_tmp564 = (w_sys_tmp565 + r_run_k_9);
	assign w_sys_tmp565 = 32'sh000013e7;
	assign w_sys_tmp570 = (w_sys_tmp571 + r_run_k_9);
	assign w_sys_tmp571 = 32'sh00001428;
	assign w_sys_tmp576 = (w_sys_tmp577 + r_run_k_9);
	assign w_sys_tmp577 = 32'sh00001448;
	assign w_sys_tmp582 = (w_sys_tmp583 + r_run_k_9);
	assign w_sys_tmp583 = 32'sh00001468;
	assign w_sys_tmp588 = (w_sys_tmp589 + r_run_k_9);
	assign w_sys_tmp589 = 32'sh000014a9;
	assign w_sys_tmp594 = (w_sys_tmp595 + r_run_k_9);
	assign w_sys_tmp595 = 32'sh000014c9;
	assign w_sys_tmp600 = (w_sys_tmp601 + r_run_k_9);
	assign w_sys_tmp601 = 32'sh000014e9;
	assign w_sys_tmp606 = (w_sys_tmp607 + r_run_k_9);
	assign w_sys_tmp607 = 32'sh0000152a;
	assign w_sys_tmp612 = (w_sys_tmp613 + r_run_k_9);
	assign w_sys_tmp613 = 32'sh0000154a;
	assign w_sys_tmp618 = (w_sys_tmp619 + r_run_k_9);
	assign w_sys_tmp619 = 32'sh0000156a;
	assign w_sys_tmp624 = (w_sys_tmp625 + r_run_k_9);
	assign w_sys_tmp625 = 32'sh000015ab;
	assign w_sys_tmp630 = (w_sys_tmp631 + r_run_k_9);
	assign w_sys_tmp631 = 32'sh000015cb;
	assign w_sys_tmp636 = (w_sys_tmp637 + r_run_k_9);
	assign w_sys_tmp637 = 32'sh000015eb;
	assign w_sys_tmp642 = (w_sys_tmp643 + r_run_k_9);
	assign w_sys_tmp643 = 32'sh0000162c;
	assign w_sys_tmp648 = (w_sys_tmp649 + r_run_k_9);
	assign w_sys_tmp649 = 32'sh0000164c;
	assign w_sys_tmp654 = (w_sys_tmp655 + r_run_k_9);
	assign w_sys_tmp655 = 32'sh0000166c;
	assign w_sys_tmp660 = (w_sys_tmp661 + r_run_k_9);
	assign w_sys_tmp661 = 32'sh000016ad;
	assign w_sys_tmp666 = (w_sys_tmp667 + r_run_k_9);
	assign w_sys_tmp667 = 32'sh000016cd;
	assign w_sys_tmp672 = (w_sys_tmp673 + r_run_k_9);
	assign w_sys_tmp673 = 32'sh000016ed;
	assign w_sys_tmp678 = (w_sys_tmp679 + r_run_k_9);
	assign w_sys_tmp679 = 32'sh0000172e;
	assign w_sys_tmp684 = (w_sys_tmp685 + r_run_k_9);
	assign w_sys_tmp685 = 32'sh0000174e;
	assign w_sys_tmp690 = (w_sys_tmp691 + r_run_k_9);
	assign w_sys_tmp691 = 32'sh0000176e;
	assign w_sys_tmp696 = (w_sys_tmp697 + r_run_k_9);
	assign w_sys_tmp697 = 32'sh000017af;
	assign w_sys_tmp702 = (w_sys_tmp703 + r_run_k_9);
	assign w_sys_tmp703 = 32'sh000017cf;
	assign w_sys_tmp708 = (w_sys_tmp709 + r_run_k_9);
	assign w_sys_tmp709 = 32'sh000017ef;
	assign w_sys_tmp714 = (w_sys_tmp715 + r_run_k_9);
	assign w_sys_tmp715 = 32'sh00001830;
	assign w_sys_tmp720 = (w_sys_tmp721 + r_run_k_9);
	assign w_sys_tmp721 = 32'sh00001850;
	assign w_sys_tmp726 = (w_sys_tmp727 + r_run_k_9);
	assign w_sys_tmp727 = 32'sh00001870;
	assign w_sys_tmp732 = (w_sys_tmp733 + r_run_k_9);
	assign w_sys_tmp733 = 32'sh000018b1;
	assign w_sys_tmp738 = (w_sys_tmp739 + r_run_k_9);
	assign w_sys_tmp739 = 32'sh000018d1;
	assign w_sys_tmp744 = (w_sys_tmp745 + r_run_k_9);
	assign w_sys_tmp745 = 32'sh000018f1;
	assign w_sys_tmp750 = (w_sys_tmp751 + r_run_k_9);
	assign w_sys_tmp751 = 32'sh00001932;
	assign w_sys_tmp756 = (w_sys_tmp757 + r_run_k_9);
	assign w_sys_tmp757 = 32'sh00001952;
	assign w_sys_tmp762 = (w_sys_tmp763 + r_run_k_9);
	assign w_sys_tmp763 = 32'sh00001972;
	assign w_sys_tmp768 = (w_sys_tmp769 + r_run_k_9);
	assign w_sys_tmp769 = 32'sh000019b3;
	assign w_sys_tmp774 = (w_sys_tmp775 + r_run_k_9);
	assign w_sys_tmp775 = 32'sh000019d3;
	assign w_sys_tmp780 = (w_sys_tmp781 + r_run_k_9);
	assign w_sys_tmp781 = 32'sh000019f3;
	assign w_sys_tmp786 = (w_sys_tmp787 + r_run_k_9);
	assign w_sys_tmp787 = 32'sh00001a34;
	assign w_sys_tmp792 = (w_sys_tmp793 + r_run_k_9);
	assign w_sys_tmp793 = 32'sh00001a54;
	assign w_sys_tmp798 = (w_sys_tmp799 + r_run_k_9);
	assign w_sys_tmp799 = 32'sh00001a74;
	assign w_sys_tmp804 = (w_sys_tmp805 + r_run_k_9);
	assign w_sys_tmp805 = 32'sh00001ab5;
	assign w_sys_tmp810 = (w_sys_tmp811 + r_run_k_9);
	assign w_sys_tmp811 = 32'sh00001ad5;
	assign w_sys_tmp816 = (w_sys_tmp817 + r_run_k_9);
	assign w_sys_tmp817 = 32'sh00001af5;
	assign w_sys_tmp822 = (w_sys_tmp823 + r_run_k_9);
	assign w_sys_tmp823 = 32'sh00001b36;
	assign w_sys_tmp828 = (w_sys_tmp829 + r_run_k_9);
	assign w_sys_tmp829 = 32'sh00001b56;
	assign w_sys_tmp834 = (w_sys_tmp835 + r_run_k_9);
	assign w_sys_tmp835 = 32'sh00001b76;
	assign w_sys_tmp840 = (w_sys_tmp841 + r_run_k_9);
	assign w_sys_tmp841 = 32'sh00001bb7;
	assign w_sys_tmp846 = (w_sys_tmp847 + r_run_k_9);
	assign w_sys_tmp847 = 32'sh00001bd7;
	assign w_sys_tmp852 = (w_sys_tmp853 + r_run_k_9);
	assign w_sys_tmp853 = 32'sh00001bf7;
	assign w_sys_tmp858 = (w_sys_tmp859 + r_run_k_9);
	assign w_sys_tmp859 = 32'sh00001c38;
	assign w_sys_tmp864 = (w_sys_tmp865 + r_run_k_9);
	assign w_sys_tmp865 = 32'sh00001c58;
	assign w_sys_tmp870 = (w_sys_tmp871 + r_run_k_9);
	assign w_sys_tmp871 = 32'sh00001c78;
	assign w_sys_tmp876 = (w_sys_tmp877 + r_run_k_9);
	assign w_sys_tmp877 = 32'sh00001cb9;
	assign w_sys_tmp882 = (w_sys_tmp883 + r_run_k_9);
	assign w_sys_tmp883 = 32'sh00001cd9;
	assign w_sys_tmp888 = (w_sys_tmp889 + r_run_k_9);
	assign w_sys_tmp889 = 32'sh00001cf9;
	assign w_sys_tmp894 = (w_sys_tmp895 + r_run_k_9);
	assign w_sys_tmp895 = 32'sh00001d3a;
	assign w_sys_tmp900 = (w_sys_tmp901 + r_run_k_9);
	assign w_sys_tmp901 = 32'sh00001d5a;
	assign w_sys_tmp906 = (w_sys_tmp907 + r_run_k_9);
	assign w_sys_tmp907 = 32'sh00001d7a;
	assign w_sys_tmp912 = (w_sys_tmp913 + r_run_k_9);
	assign w_sys_tmp913 = 32'sh00001dbb;
	assign w_sys_tmp918 = (w_sys_tmp919 + r_run_k_9);
	assign w_sys_tmp919 = 32'sh00001ddb;
	assign w_sys_tmp924 = (w_sys_tmp925 + r_run_k_9);
	assign w_sys_tmp925 = 32'sh00001dfb;
	assign w_sys_tmp930 = (w_sys_tmp931 + r_run_k_9);
	assign w_sys_tmp931 = 32'sh00001e3c;
	assign w_sys_tmp936 = (w_sys_tmp937 + r_run_k_9);
	assign w_sys_tmp937 = 32'sh00001e5c;
	assign w_sys_tmp942 = (w_sys_tmp943 + r_run_k_9);
	assign w_sys_tmp943 = 32'sh00001e7c;
	assign w_sys_tmp948 = (w_sys_tmp949 + r_run_k_9);
	assign w_sys_tmp949 = 32'sh00001ebd;
	assign w_sys_tmp954 = (w_sys_tmp955 + r_run_k_9);
	assign w_sys_tmp955 = 32'sh00001edd;
	assign w_sys_tmp960 = (w_sys_tmp961 + r_run_k_9);
	assign w_sys_tmp961 = 32'sh00001efd;
	assign w_sys_tmp966 = (w_sys_tmp967 + r_run_k_9);
	assign w_sys_tmp967 = 32'sh00001f3e;
	assign w_sys_tmp972 = (w_sys_tmp973 + r_run_k_9);
	assign w_sys_tmp973 = 32'sh00001f5e;
	assign w_sys_tmp978 = (w_sys_tmp979 + r_run_k_9);
	assign w_sys_tmp979 = 32'sh00001f7e;
	assign w_sys_tmp984 = (w_sys_tmp985 + r_run_k_9);
	assign w_sys_tmp985 = 32'sh00001fbf;
	assign w_sys_tmp990 = (w_sys_tmp991 + r_run_k_9);
	assign w_sys_tmp991 = 32'sh00001fdf;
	assign w_sys_tmp996 = (w_sys_tmp997 + r_run_k_9);
	assign w_sys_tmp997 = 32'sh00001fff;
	assign w_sys_tmp1002 = (w_sys_tmp1003 + r_run_k_9);
	assign w_sys_tmp1003 = 32'sh00002040;
	assign w_sys_tmp1008 = (w_sys_tmp1009 + r_run_k_9);
	assign w_sys_tmp1009 = 32'sh00002060;
	assign w_sys_tmp1014 = (w_sys_tmp1015 + r_run_k_9);
	assign w_sys_tmp1015 = 32'sh00002080;
	assign w_sys_tmp1020 = (w_sys_tmp1021 + r_run_k_9);
	assign w_sys_tmp1021 = 32'sh000020c1;
	assign w_sys_tmp1026 = (w_sys_tmp1027 + r_run_k_9);
	assign w_sys_tmp1027 = 32'sh000020e1;
	assign w_sys_tmp1032 = (w_sys_tmp1033 + r_run_k_9);
	assign w_sys_tmp1033 = 32'sh00002101;
	assign w_sys_tmp1037 = (r_run_k_9 + w_sys_intOne);
	assign w_sys_tmp1038 = 32'sh00000040;
	assign w_sys_tmp1039 = ( !w_sys_tmp1040 );
	assign w_sys_tmp1040 = (w_sys_tmp1041 < r_run_k_9);
	assign w_sys_tmp1041 = 32'sh00000081;
	assign w_sys_tmp1044 = (w_sys_tmp1045 + r_run_k_9);
	assign w_sys_tmp1045 = 32'sh00000081;
	assign w_sys_tmp1046 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1050 = (w_sys_tmp1051 + r_run_k_9);
	assign w_sys_tmp1051 = 32'sh00000102;
	assign w_sys_tmp1056 = (w_sys_tmp1057 + r_run_k_9);
	assign w_sys_tmp1057 = 32'sh00000183;
	assign w_sys_tmp1062 = (w_sys_tmp1063 + r_run_k_9);
	assign w_sys_tmp1063 = 32'sh00000204;
	assign w_sys_tmp1068 = (w_sys_tmp1069 + r_run_k_9);
	assign w_sys_tmp1069 = 32'sh00000285;
	assign w_sys_tmp1074 = (w_sys_tmp1075 + r_run_k_9);
	assign w_sys_tmp1075 = 32'sh00000306;
	assign w_sys_tmp1080 = (w_sys_tmp1081 + r_run_k_9);
	assign w_sys_tmp1081 = 32'sh00000387;
	assign w_sys_tmp1086 = (w_sys_tmp1087 + r_run_k_9);
	assign w_sys_tmp1087 = 32'sh00000408;
	assign w_sys_tmp1092 = (w_sys_tmp1093 + r_run_k_9);
	assign w_sys_tmp1093 = 32'sh00000489;
	assign w_sys_tmp1098 = (w_sys_tmp1099 + r_run_k_9);
	assign w_sys_tmp1099 = 32'sh0000050a;
	assign w_sys_tmp1104 = (w_sys_tmp1105 + r_run_k_9);
	assign w_sys_tmp1105 = 32'sh0000058b;
	assign w_sys_tmp1110 = (w_sys_tmp1111 + r_run_k_9);
	assign w_sys_tmp1111 = 32'sh0000060c;
	assign w_sys_tmp1116 = (w_sys_tmp1117 + r_run_k_9);
	assign w_sys_tmp1117 = 32'sh0000068d;
	assign w_sys_tmp1122 = (w_sys_tmp1123 + r_run_k_9);
	assign w_sys_tmp1123 = 32'sh0000070e;
	assign w_sys_tmp1128 = (w_sys_tmp1129 + r_run_k_9);
	assign w_sys_tmp1129 = 32'sh0000078f;
	assign w_sys_tmp1134 = (w_sys_tmp1135 + r_run_k_9);
	assign w_sys_tmp1135 = 32'sh00000810;
	assign w_sys_tmp1140 = (w_sys_tmp1141 + r_run_k_9);
	assign w_sys_tmp1141 = 32'sh00000891;
	assign w_sys_tmp1146 = (w_sys_tmp1147 + r_run_k_9);
	assign w_sys_tmp1147 = 32'sh00000912;
	assign w_sys_tmp1152 = (w_sys_tmp1153 + r_run_k_9);
	assign w_sys_tmp1153 = 32'sh00000993;
	assign w_sys_tmp1158 = (w_sys_tmp1159 + r_run_k_9);
	assign w_sys_tmp1159 = 32'sh00000a14;
	assign w_sys_tmp1164 = (w_sys_tmp1165 + r_run_k_9);
	assign w_sys_tmp1165 = 32'sh00000a95;
	assign w_sys_tmp1170 = (w_sys_tmp1171 + r_run_k_9);
	assign w_sys_tmp1171 = 32'sh00000b16;
	assign w_sys_tmp1176 = (w_sys_tmp1177 + r_run_k_9);
	assign w_sys_tmp1177 = 32'sh00000b97;
	assign w_sys_tmp1182 = (w_sys_tmp1183 + r_run_k_9);
	assign w_sys_tmp1183 = 32'sh00000c18;
	assign w_sys_tmp1188 = (w_sys_tmp1189 + r_run_k_9);
	assign w_sys_tmp1189 = 32'sh00000c99;
	assign w_sys_tmp1194 = (w_sys_tmp1195 + r_run_k_9);
	assign w_sys_tmp1195 = 32'sh00000d1a;
	assign w_sys_tmp1200 = (w_sys_tmp1201 + r_run_k_9);
	assign w_sys_tmp1201 = 32'sh00000d9b;
	assign w_sys_tmp1206 = (w_sys_tmp1207 + r_run_k_9);
	assign w_sys_tmp1207 = 32'sh00000e1c;
	assign w_sys_tmp1212 = (w_sys_tmp1213 + r_run_k_9);
	assign w_sys_tmp1213 = 32'sh00000e9d;
	assign w_sys_tmp1218 = (w_sys_tmp1219 + r_run_k_9);
	assign w_sys_tmp1219 = 32'sh00000f1e;
	assign w_sys_tmp1224 = (w_sys_tmp1225 + r_run_k_9);
	assign w_sys_tmp1225 = 32'sh00000f9f;
	assign w_sys_tmp1230 = (w_sys_tmp1231 + r_run_k_9);
	assign w_sys_tmp1231 = 32'sh00001020;
	assign w_sys_tmp1236 = (w_sys_tmp1237 + r_run_k_9);
	assign w_sys_tmp1237 = 32'sh000010a1;
	assign w_sys_tmp1248 = (w_sys_tmp1249 + r_run_k_9);
	assign w_sys_tmp1249 = 32'sh00001040;
	assign w_sys_tmp1254 = (w_sys_tmp1255 + r_run_k_9);
	assign w_sys_tmp1255 = 32'sh00001060;
	assign w_sys_tmp1266 = (w_sys_tmp1267 + r_run_k_9);
	assign w_sys_tmp1267 = 32'sh000010c1;
	assign w_sys_tmp1272 = (w_sys_tmp1273 + r_run_k_9);
	assign w_sys_tmp1273 = 32'sh000010e1;
	assign w_sys_tmp1278 = (w_sys_tmp1279 + r_run_k_9);
	assign w_sys_tmp1279 = 32'sh00001122;
	assign w_sys_tmp1284 = (w_sys_tmp1285 + r_run_k_9);
	assign w_sys_tmp1285 = 32'sh00001142;
	assign w_sys_tmp1290 = (w_sys_tmp1291 + r_run_k_9);
	assign w_sys_tmp1291 = 32'sh00001162;
	assign w_sys_tmp1296 = (w_sys_tmp1297 + r_run_k_9);
	assign w_sys_tmp1297 = 32'sh000011a3;
	assign w_sys_tmp1302 = (w_sys_tmp1303 + r_run_k_9);
	assign w_sys_tmp1303 = 32'sh000011c3;
	assign w_sys_tmp1308 = (w_sys_tmp1309 + r_run_k_9);
	assign w_sys_tmp1309 = 32'sh000011e3;
	assign w_sys_tmp1314 = (w_sys_tmp1315 + r_run_k_9);
	assign w_sys_tmp1315 = 32'sh00001224;
	assign w_sys_tmp1320 = (w_sys_tmp1321 + r_run_k_9);
	assign w_sys_tmp1321 = 32'sh00001244;
	assign w_sys_tmp1326 = (w_sys_tmp1327 + r_run_k_9);
	assign w_sys_tmp1327 = 32'sh00001264;
	assign w_sys_tmp1332 = (w_sys_tmp1333 + r_run_k_9);
	assign w_sys_tmp1333 = 32'sh000012a5;
	assign w_sys_tmp1338 = (w_sys_tmp1339 + r_run_k_9);
	assign w_sys_tmp1339 = 32'sh000012c5;
	assign w_sys_tmp1344 = (w_sys_tmp1345 + r_run_k_9);
	assign w_sys_tmp1345 = 32'sh000012e5;
	assign w_sys_tmp1350 = (w_sys_tmp1351 + r_run_k_9);
	assign w_sys_tmp1351 = 32'sh00001326;
	assign w_sys_tmp1356 = (w_sys_tmp1357 + r_run_k_9);
	assign w_sys_tmp1357 = 32'sh00001346;
	assign w_sys_tmp1362 = (w_sys_tmp1363 + r_run_k_9);
	assign w_sys_tmp1363 = 32'sh00001366;
	assign w_sys_tmp1368 = (w_sys_tmp1369 + r_run_k_9);
	assign w_sys_tmp1369 = 32'sh000013a7;
	assign w_sys_tmp1374 = (w_sys_tmp1375 + r_run_k_9);
	assign w_sys_tmp1375 = 32'sh000013c7;
	assign w_sys_tmp1380 = (w_sys_tmp1381 + r_run_k_9);
	assign w_sys_tmp1381 = 32'sh000013e7;
	assign w_sys_tmp1386 = (w_sys_tmp1387 + r_run_k_9);
	assign w_sys_tmp1387 = 32'sh00001428;
	assign w_sys_tmp1392 = (w_sys_tmp1393 + r_run_k_9);
	assign w_sys_tmp1393 = 32'sh00001448;
	assign w_sys_tmp1398 = (w_sys_tmp1399 + r_run_k_9);
	assign w_sys_tmp1399 = 32'sh00001468;
	assign w_sys_tmp1404 = (w_sys_tmp1405 + r_run_k_9);
	assign w_sys_tmp1405 = 32'sh000014a9;
	assign w_sys_tmp1410 = (w_sys_tmp1411 + r_run_k_9);
	assign w_sys_tmp1411 = 32'sh000014c9;
	assign w_sys_tmp1416 = (w_sys_tmp1417 + r_run_k_9);
	assign w_sys_tmp1417 = 32'sh000014e9;
	assign w_sys_tmp1422 = (w_sys_tmp1423 + r_run_k_9);
	assign w_sys_tmp1423 = 32'sh0000152a;
	assign w_sys_tmp1428 = (w_sys_tmp1429 + r_run_k_9);
	assign w_sys_tmp1429 = 32'sh0000154a;
	assign w_sys_tmp1434 = (w_sys_tmp1435 + r_run_k_9);
	assign w_sys_tmp1435 = 32'sh0000156a;
	assign w_sys_tmp1440 = (w_sys_tmp1441 + r_run_k_9);
	assign w_sys_tmp1441 = 32'sh000015ab;
	assign w_sys_tmp1446 = (w_sys_tmp1447 + r_run_k_9);
	assign w_sys_tmp1447 = 32'sh000015cb;
	assign w_sys_tmp1452 = (w_sys_tmp1453 + r_run_k_9);
	assign w_sys_tmp1453 = 32'sh000015eb;
	assign w_sys_tmp1458 = (w_sys_tmp1459 + r_run_k_9);
	assign w_sys_tmp1459 = 32'sh0000162c;
	assign w_sys_tmp1464 = (w_sys_tmp1465 + r_run_k_9);
	assign w_sys_tmp1465 = 32'sh0000164c;
	assign w_sys_tmp1470 = (w_sys_tmp1471 + r_run_k_9);
	assign w_sys_tmp1471 = 32'sh0000166c;
	assign w_sys_tmp1476 = (w_sys_tmp1477 + r_run_k_9);
	assign w_sys_tmp1477 = 32'sh000016ad;
	assign w_sys_tmp1482 = (w_sys_tmp1483 + r_run_k_9);
	assign w_sys_tmp1483 = 32'sh000016cd;
	assign w_sys_tmp1488 = (w_sys_tmp1489 + r_run_k_9);
	assign w_sys_tmp1489 = 32'sh000016ed;
	assign w_sys_tmp1494 = (w_sys_tmp1495 + r_run_k_9);
	assign w_sys_tmp1495 = 32'sh0000172e;
	assign w_sys_tmp1500 = (w_sys_tmp1501 + r_run_k_9);
	assign w_sys_tmp1501 = 32'sh0000174e;
	assign w_sys_tmp1506 = (w_sys_tmp1507 + r_run_k_9);
	assign w_sys_tmp1507 = 32'sh0000176e;
	assign w_sys_tmp1512 = (w_sys_tmp1513 + r_run_k_9);
	assign w_sys_tmp1513 = 32'sh000017af;
	assign w_sys_tmp1518 = (w_sys_tmp1519 + r_run_k_9);
	assign w_sys_tmp1519 = 32'sh000017cf;
	assign w_sys_tmp1524 = (w_sys_tmp1525 + r_run_k_9);
	assign w_sys_tmp1525 = 32'sh000017ef;
	assign w_sys_tmp1530 = (w_sys_tmp1531 + r_run_k_9);
	assign w_sys_tmp1531 = 32'sh00001830;
	assign w_sys_tmp1536 = (w_sys_tmp1537 + r_run_k_9);
	assign w_sys_tmp1537 = 32'sh00001850;
	assign w_sys_tmp1542 = (w_sys_tmp1543 + r_run_k_9);
	assign w_sys_tmp1543 = 32'sh00001870;
	assign w_sys_tmp1548 = (w_sys_tmp1549 + r_run_k_9);
	assign w_sys_tmp1549 = 32'sh000018b1;
	assign w_sys_tmp1554 = (w_sys_tmp1555 + r_run_k_9);
	assign w_sys_tmp1555 = 32'sh000018d1;
	assign w_sys_tmp1560 = (w_sys_tmp1561 + r_run_k_9);
	assign w_sys_tmp1561 = 32'sh000018f1;
	assign w_sys_tmp1566 = (w_sys_tmp1567 + r_run_k_9);
	assign w_sys_tmp1567 = 32'sh00001932;
	assign w_sys_tmp1572 = (w_sys_tmp1573 + r_run_k_9);
	assign w_sys_tmp1573 = 32'sh00001952;
	assign w_sys_tmp1578 = (w_sys_tmp1579 + r_run_k_9);
	assign w_sys_tmp1579 = 32'sh00001972;
	assign w_sys_tmp1584 = (w_sys_tmp1585 + r_run_k_9);
	assign w_sys_tmp1585 = 32'sh000019b3;
	assign w_sys_tmp1590 = (w_sys_tmp1591 + r_run_k_9);
	assign w_sys_tmp1591 = 32'sh000019d3;
	assign w_sys_tmp1596 = (w_sys_tmp1597 + r_run_k_9);
	assign w_sys_tmp1597 = 32'sh000019f3;
	assign w_sys_tmp1602 = (w_sys_tmp1603 + r_run_k_9);
	assign w_sys_tmp1603 = 32'sh00001a34;
	assign w_sys_tmp1608 = (w_sys_tmp1609 + r_run_k_9);
	assign w_sys_tmp1609 = 32'sh00001a54;
	assign w_sys_tmp1614 = (w_sys_tmp1615 + r_run_k_9);
	assign w_sys_tmp1615 = 32'sh00001a74;
	assign w_sys_tmp1620 = (w_sys_tmp1621 + r_run_k_9);
	assign w_sys_tmp1621 = 32'sh00001ab5;
	assign w_sys_tmp1626 = (w_sys_tmp1627 + r_run_k_9);
	assign w_sys_tmp1627 = 32'sh00001ad5;
	assign w_sys_tmp1632 = (w_sys_tmp1633 + r_run_k_9);
	assign w_sys_tmp1633 = 32'sh00001af5;
	assign w_sys_tmp1638 = (w_sys_tmp1639 + r_run_k_9);
	assign w_sys_tmp1639 = 32'sh00001b36;
	assign w_sys_tmp1644 = (w_sys_tmp1645 + r_run_k_9);
	assign w_sys_tmp1645 = 32'sh00001b56;
	assign w_sys_tmp1650 = (w_sys_tmp1651 + r_run_k_9);
	assign w_sys_tmp1651 = 32'sh00001b76;
	assign w_sys_tmp1656 = (w_sys_tmp1657 + r_run_k_9);
	assign w_sys_tmp1657 = 32'sh00001bb7;
	assign w_sys_tmp1662 = (w_sys_tmp1663 + r_run_k_9);
	assign w_sys_tmp1663 = 32'sh00001bd7;
	assign w_sys_tmp1668 = (w_sys_tmp1669 + r_run_k_9);
	assign w_sys_tmp1669 = 32'sh00001bf7;
	assign w_sys_tmp1674 = (w_sys_tmp1675 + r_run_k_9);
	assign w_sys_tmp1675 = 32'sh00001c38;
	assign w_sys_tmp1680 = (w_sys_tmp1681 + r_run_k_9);
	assign w_sys_tmp1681 = 32'sh00001c58;
	assign w_sys_tmp1686 = (w_sys_tmp1687 + r_run_k_9);
	assign w_sys_tmp1687 = 32'sh00001c78;
	assign w_sys_tmp1692 = (w_sys_tmp1693 + r_run_k_9);
	assign w_sys_tmp1693 = 32'sh00001cb9;
	assign w_sys_tmp1698 = (w_sys_tmp1699 + r_run_k_9);
	assign w_sys_tmp1699 = 32'sh00001cd9;
	assign w_sys_tmp1704 = (w_sys_tmp1705 + r_run_k_9);
	assign w_sys_tmp1705 = 32'sh00001cf9;
	assign w_sys_tmp1710 = (w_sys_tmp1711 + r_run_k_9);
	assign w_sys_tmp1711 = 32'sh00001d3a;
	assign w_sys_tmp1716 = (w_sys_tmp1717 + r_run_k_9);
	assign w_sys_tmp1717 = 32'sh00001d5a;
	assign w_sys_tmp1722 = (w_sys_tmp1723 + r_run_k_9);
	assign w_sys_tmp1723 = 32'sh00001d7a;
	assign w_sys_tmp1728 = (w_sys_tmp1729 + r_run_k_9);
	assign w_sys_tmp1729 = 32'sh00001dbb;
	assign w_sys_tmp1734 = (w_sys_tmp1735 + r_run_k_9);
	assign w_sys_tmp1735 = 32'sh00001ddb;
	assign w_sys_tmp1740 = (w_sys_tmp1741 + r_run_k_9);
	assign w_sys_tmp1741 = 32'sh00001dfb;
	assign w_sys_tmp1746 = (w_sys_tmp1747 + r_run_k_9);
	assign w_sys_tmp1747 = 32'sh00001e3c;
	assign w_sys_tmp1752 = (w_sys_tmp1753 + r_run_k_9);
	assign w_sys_tmp1753 = 32'sh00001e5c;
	assign w_sys_tmp1758 = (w_sys_tmp1759 + r_run_k_9);
	assign w_sys_tmp1759 = 32'sh00001e7c;
	assign w_sys_tmp1764 = (w_sys_tmp1765 + r_run_k_9);
	assign w_sys_tmp1765 = 32'sh00001ebd;
	assign w_sys_tmp1770 = (w_sys_tmp1771 + r_run_k_9);
	assign w_sys_tmp1771 = 32'sh00001edd;
	assign w_sys_tmp1776 = (w_sys_tmp1777 + r_run_k_9);
	assign w_sys_tmp1777 = 32'sh00001efd;
	assign w_sys_tmp1782 = (w_sys_tmp1783 + r_run_k_9);
	assign w_sys_tmp1783 = 32'sh00001f3e;
	assign w_sys_tmp1788 = (w_sys_tmp1789 + r_run_k_9);
	assign w_sys_tmp1789 = 32'sh00001f5e;
	assign w_sys_tmp1794 = (w_sys_tmp1795 + r_run_k_9);
	assign w_sys_tmp1795 = 32'sh00001f7e;
	assign w_sys_tmp1800 = (w_sys_tmp1801 + r_run_k_9);
	assign w_sys_tmp1801 = 32'sh00001fbf;
	assign w_sys_tmp1806 = (w_sys_tmp1807 + r_run_k_9);
	assign w_sys_tmp1807 = 32'sh00001fdf;
	assign w_sys_tmp1812 = (w_sys_tmp1813 + r_run_k_9);
	assign w_sys_tmp1813 = 32'sh00001fff;
	assign w_sys_tmp1818 = (w_sys_tmp1819 + r_run_k_9);
	assign w_sys_tmp1819 = 32'sh00002040;
	assign w_sys_tmp1824 = (w_sys_tmp1825 + r_run_k_9);
	assign w_sys_tmp1825 = 32'sh00002060;
	assign w_sys_tmp1830 = (w_sys_tmp1831 + r_run_k_9);
	assign w_sys_tmp1831 = 32'sh00002080;
	assign w_sys_tmp1836 = (w_sys_tmp1837 + r_run_k_9);
	assign w_sys_tmp1837 = 32'sh000020c1;
	assign w_sys_tmp1842 = (w_sys_tmp1843 + r_run_k_9);
	assign w_sys_tmp1843 = 32'sh000020e1;
	assign w_sys_tmp1848 = (w_sys_tmp1849 + r_run_k_9);
	assign w_sys_tmp1849 = 32'sh00002101;
	assign w_sys_tmp1853 = (r_run_k_9 + w_sys_intOne);
	assign w_sys_tmp1854 = 32'sh00000002;
	assign w_sys_tmp1855 = ( !w_sys_tmp1856 );
	assign w_sys_tmp1856 = (w_sys_tmp1857 < r_run_k_9);
	assign w_sys_tmp1857 = 32'sh00000040;
	assign w_sys_tmp1860 = (w_sys_tmp1861 + r_run_k_9);
	assign w_sys_tmp1861 = 32'sh00000102;
	assign w_sys_tmp1862 = w_sub00_result_dataout;
	assign w_sys_tmp1866 = (w_sys_tmp1867 + r_run_k_9);
	assign w_sys_tmp1867 = 32'sh00000183;
	assign w_sys_tmp1872 = (w_sys_tmp1873 + r_run_k_9);
	assign w_sys_tmp1873 = 32'sh00000204;
	assign w_sys_tmp1878 = (w_sys_tmp1879 + r_run_k_9);
	assign w_sys_tmp1879 = 32'sh00000285;
	assign w_sys_tmp1884 = (w_sys_tmp1885 + r_run_k_9);
	assign w_sys_tmp1885 = 32'sh00000306;
	assign w_sys_tmp1890 = (w_sys_tmp1891 + r_run_k_9);
	assign w_sys_tmp1891 = 32'sh00000387;
	assign w_sys_tmp1896 = (w_sys_tmp1897 + r_run_k_9);
	assign w_sys_tmp1897 = 32'sh00000408;
	assign w_sys_tmp1902 = (w_sys_tmp1903 + r_run_k_9);
	assign w_sys_tmp1903 = 32'sh00000489;
	assign w_sys_tmp1908 = (w_sys_tmp1909 + r_run_k_9);
	assign w_sys_tmp1909 = 32'sh0000050a;
	assign w_sys_tmp1914 = (w_sys_tmp1915 + r_run_k_9);
	assign w_sys_tmp1915 = 32'sh0000058b;
	assign w_sys_tmp1920 = (w_sys_tmp1921 + r_run_k_9);
	assign w_sys_tmp1921 = 32'sh0000060c;
	assign w_sys_tmp1926 = (w_sys_tmp1927 + r_run_k_9);
	assign w_sys_tmp1927 = 32'sh0000068d;
	assign w_sys_tmp1932 = (w_sys_tmp1933 + r_run_k_9);
	assign w_sys_tmp1933 = 32'sh0000070e;
	assign w_sys_tmp1938 = (w_sys_tmp1939 + r_run_k_9);
	assign w_sys_tmp1939 = 32'sh0000078f;
	assign w_sys_tmp1944 = (w_sys_tmp1945 + r_run_k_9);
	assign w_sys_tmp1945 = 32'sh00000810;
	assign w_sys_tmp1950 = (w_sys_tmp1951 + r_run_k_9);
	assign w_sys_tmp1951 = 32'sh00000891;
	assign w_sys_tmp1956 = (w_sys_tmp1957 + r_run_k_9);
	assign w_sys_tmp1957 = 32'sh00000912;
	assign w_sys_tmp1962 = (w_sys_tmp1963 + r_run_k_9);
	assign w_sys_tmp1963 = 32'sh00000993;
	assign w_sys_tmp1968 = (w_sys_tmp1969 + r_run_k_9);
	assign w_sys_tmp1969 = 32'sh00000a14;
	assign w_sys_tmp1974 = (w_sys_tmp1975 + r_run_k_9);
	assign w_sys_tmp1975 = 32'sh00000a95;
	assign w_sys_tmp1980 = (w_sys_tmp1981 + r_run_k_9);
	assign w_sys_tmp1981 = 32'sh00000b16;
	assign w_sys_tmp1986 = (w_sys_tmp1987 + r_run_k_9);
	assign w_sys_tmp1987 = 32'sh00000b97;
	assign w_sys_tmp1992 = (w_sys_tmp1993 + r_run_k_9);
	assign w_sys_tmp1993 = 32'sh00000c18;
	assign w_sys_tmp1998 = (w_sys_tmp1999 + r_run_k_9);
	assign w_sys_tmp1999 = 32'sh00000c99;
	assign w_sys_tmp2004 = (w_sys_tmp2005 + r_run_k_9);
	assign w_sys_tmp2005 = 32'sh00000d1a;
	assign w_sys_tmp2010 = (w_sys_tmp2011 + r_run_k_9);
	assign w_sys_tmp2011 = 32'sh00000d9b;
	assign w_sys_tmp2016 = (w_sys_tmp2017 + r_run_k_9);
	assign w_sys_tmp2017 = 32'sh00000e1c;
	assign w_sys_tmp2022 = (w_sys_tmp2023 + r_run_k_9);
	assign w_sys_tmp2023 = 32'sh00000e9d;
	assign w_sys_tmp2028 = (w_sys_tmp2029 + r_run_k_9);
	assign w_sys_tmp2029 = 32'sh00000f1e;
	assign w_sys_tmp2034 = (w_sys_tmp2035 + r_run_k_9);
	assign w_sys_tmp2035 = 32'sh00000f9f;
	assign w_sys_tmp2040 = (w_sys_tmp2041 + r_run_k_9);
	assign w_sys_tmp2041 = 32'sh00001020;
	assign w_sys_tmp2046 = (w_sys_tmp2047 + r_run_k_9);
	assign w_sys_tmp2047 = 32'sh000010a1;
	assign w_sys_tmp2051 = (w_sys_tmp2052 + r_run_k_9);
	assign w_sys_tmp2052 = 32'sh000010c1;
	assign w_sys_tmp2056 = (w_sys_tmp2057 + r_run_k_9);
	assign w_sys_tmp2057 = 32'sh000010e1;
	assign w_sys_tmp2061 = (w_sys_tmp2062 + r_run_k_9);
	assign w_sys_tmp2062 = 32'sh00001122;
	assign w_sys_tmp2066 = (w_sys_tmp2067 + r_run_k_9);
	assign w_sys_tmp2067 = 32'sh00001142;
	assign w_sys_tmp2071 = (w_sys_tmp2072 + r_run_k_9);
	assign w_sys_tmp2072 = 32'sh00001162;
	assign w_sys_tmp2076 = (w_sys_tmp2077 + r_run_k_9);
	assign w_sys_tmp2077 = 32'sh000011a3;
	assign w_sys_tmp2081 = (w_sys_tmp2082 + r_run_k_9);
	assign w_sys_tmp2082 = 32'sh000011c3;
	assign w_sys_tmp2086 = (w_sys_tmp2087 + r_run_k_9);
	assign w_sys_tmp2087 = 32'sh000011e3;
	assign w_sys_tmp2091 = (w_sys_tmp2092 + r_run_k_9);
	assign w_sys_tmp2092 = 32'sh00001224;
	assign w_sys_tmp2096 = (w_sys_tmp2097 + r_run_k_9);
	assign w_sys_tmp2097 = 32'sh00001244;
	assign w_sys_tmp2101 = (w_sys_tmp2102 + r_run_k_9);
	assign w_sys_tmp2102 = 32'sh00001264;
	assign w_sys_tmp2106 = (w_sys_tmp2107 + r_run_k_9);
	assign w_sys_tmp2107 = 32'sh000012a5;
	assign w_sys_tmp2111 = (w_sys_tmp2112 + r_run_k_9);
	assign w_sys_tmp2112 = 32'sh000012c5;
	assign w_sys_tmp2116 = (w_sys_tmp2117 + r_run_k_9);
	assign w_sys_tmp2117 = 32'sh000012e5;
	assign w_sys_tmp2121 = (w_sys_tmp2122 + r_run_k_9);
	assign w_sys_tmp2122 = 32'sh00001326;
	assign w_sys_tmp2126 = (w_sys_tmp2127 + r_run_k_9);
	assign w_sys_tmp2127 = 32'sh00001346;
	assign w_sys_tmp2131 = (w_sys_tmp2132 + r_run_k_9);
	assign w_sys_tmp2132 = 32'sh00001366;
	assign w_sys_tmp2136 = (w_sys_tmp2137 + r_run_k_9);
	assign w_sys_tmp2137 = 32'sh000013a7;
	assign w_sys_tmp2141 = (w_sys_tmp2142 + r_run_k_9);
	assign w_sys_tmp2142 = 32'sh000013c7;
	assign w_sys_tmp2146 = (w_sys_tmp2147 + r_run_k_9);
	assign w_sys_tmp2147 = 32'sh000013e7;
	assign w_sys_tmp2151 = (w_sys_tmp2152 + r_run_k_9);
	assign w_sys_tmp2152 = 32'sh00001428;
	assign w_sys_tmp2156 = (w_sys_tmp2157 + r_run_k_9);
	assign w_sys_tmp2157 = 32'sh00001448;
	assign w_sys_tmp2161 = (w_sys_tmp2162 + r_run_k_9);
	assign w_sys_tmp2162 = 32'sh00001468;
	assign w_sys_tmp2166 = (w_sys_tmp2167 + r_run_k_9);
	assign w_sys_tmp2167 = 32'sh000014a9;
	assign w_sys_tmp2171 = (w_sys_tmp2172 + r_run_k_9);
	assign w_sys_tmp2172 = 32'sh000014c9;
	assign w_sys_tmp2176 = (w_sys_tmp2177 + r_run_k_9);
	assign w_sys_tmp2177 = 32'sh000014e9;
	assign w_sys_tmp2181 = (w_sys_tmp2182 + r_run_k_9);
	assign w_sys_tmp2182 = 32'sh0000152a;
	assign w_sys_tmp2186 = (w_sys_tmp2187 + r_run_k_9);
	assign w_sys_tmp2187 = 32'sh0000154a;
	assign w_sys_tmp2191 = (w_sys_tmp2192 + r_run_k_9);
	assign w_sys_tmp2192 = 32'sh0000156a;
	assign w_sys_tmp2196 = (w_sys_tmp2197 + r_run_k_9);
	assign w_sys_tmp2197 = 32'sh000015ab;
	assign w_sys_tmp2201 = (w_sys_tmp2202 + r_run_k_9);
	assign w_sys_tmp2202 = 32'sh000015cb;
	assign w_sys_tmp2206 = (w_sys_tmp2207 + r_run_k_9);
	assign w_sys_tmp2207 = 32'sh000015eb;
	assign w_sys_tmp2211 = (w_sys_tmp2212 + r_run_k_9);
	assign w_sys_tmp2212 = 32'sh0000162c;
	assign w_sys_tmp2216 = (w_sys_tmp2217 + r_run_k_9);
	assign w_sys_tmp2217 = 32'sh0000164c;
	assign w_sys_tmp2221 = (w_sys_tmp2222 + r_run_k_9);
	assign w_sys_tmp2222 = 32'sh0000166c;
	assign w_sys_tmp2226 = (w_sys_tmp2227 + r_run_k_9);
	assign w_sys_tmp2227 = 32'sh000016ad;
	assign w_sys_tmp2231 = (w_sys_tmp2232 + r_run_k_9);
	assign w_sys_tmp2232 = 32'sh000016cd;
	assign w_sys_tmp2236 = (w_sys_tmp2237 + r_run_k_9);
	assign w_sys_tmp2237 = 32'sh000016ed;
	assign w_sys_tmp2241 = (w_sys_tmp2242 + r_run_k_9);
	assign w_sys_tmp2242 = 32'sh0000172e;
	assign w_sys_tmp2246 = (w_sys_tmp2247 + r_run_k_9);
	assign w_sys_tmp2247 = 32'sh0000174e;
	assign w_sys_tmp2251 = (w_sys_tmp2252 + r_run_k_9);
	assign w_sys_tmp2252 = 32'sh0000176e;
	assign w_sys_tmp2256 = (w_sys_tmp2257 + r_run_k_9);
	assign w_sys_tmp2257 = 32'sh000017af;
	assign w_sys_tmp2261 = (w_sys_tmp2262 + r_run_k_9);
	assign w_sys_tmp2262 = 32'sh000017cf;
	assign w_sys_tmp2266 = (w_sys_tmp2267 + r_run_k_9);
	assign w_sys_tmp2267 = 32'sh000017ef;
	assign w_sys_tmp2271 = (w_sys_tmp2272 + r_run_k_9);
	assign w_sys_tmp2272 = 32'sh00001830;
	assign w_sys_tmp2276 = (w_sys_tmp2277 + r_run_k_9);
	assign w_sys_tmp2277 = 32'sh00001850;
	assign w_sys_tmp2281 = (w_sys_tmp2282 + r_run_k_9);
	assign w_sys_tmp2282 = 32'sh00001870;
	assign w_sys_tmp2286 = (w_sys_tmp2287 + r_run_k_9);
	assign w_sys_tmp2287 = 32'sh000018b1;
	assign w_sys_tmp2291 = (w_sys_tmp2292 + r_run_k_9);
	assign w_sys_tmp2292 = 32'sh000018d1;
	assign w_sys_tmp2296 = (w_sys_tmp2297 + r_run_k_9);
	assign w_sys_tmp2297 = 32'sh000018f1;
	assign w_sys_tmp2301 = (w_sys_tmp2302 + r_run_k_9);
	assign w_sys_tmp2302 = 32'sh00001932;
	assign w_sys_tmp2306 = (w_sys_tmp2307 + r_run_k_9);
	assign w_sys_tmp2307 = 32'sh00001952;
	assign w_sys_tmp2311 = (w_sys_tmp2312 + r_run_k_9);
	assign w_sys_tmp2312 = 32'sh00001972;
	assign w_sys_tmp2316 = (w_sys_tmp2317 + r_run_k_9);
	assign w_sys_tmp2317 = 32'sh000019b3;
	assign w_sys_tmp2321 = (w_sys_tmp2322 + r_run_k_9);
	assign w_sys_tmp2322 = 32'sh000019d3;
	assign w_sys_tmp2326 = (w_sys_tmp2327 + r_run_k_9);
	assign w_sys_tmp2327 = 32'sh000019f3;
	assign w_sys_tmp2331 = (w_sys_tmp2332 + r_run_k_9);
	assign w_sys_tmp2332 = 32'sh00001a34;
	assign w_sys_tmp2336 = (w_sys_tmp2337 + r_run_k_9);
	assign w_sys_tmp2337 = 32'sh00001a54;
	assign w_sys_tmp2341 = (w_sys_tmp2342 + r_run_k_9);
	assign w_sys_tmp2342 = 32'sh00001a74;
	assign w_sys_tmp2346 = (w_sys_tmp2347 + r_run_k_9);
	assign w_sys_tmp2347 = 32'sh00001ab5;
	assign w_sys_tmp2351 = (w_sys_tmp2352 + r_run_k_9);
	assign w_sys_tmp2352 = 32'sh00001ad5;
	assign w_sys_tmp2356 = (w_sys_tmp2357 + r_run_k_9);
	assign w_sys_tmp2357 = 32'sh00001af5;
	assign w_sys_tmp2361 = (w_sys_tmp2362 + r_run_k_9);
	assign w_sys_tmp2362 = 32'sh00001b36;
	assign w_sys_tmp2366 = (w_sys_tmp2367 + r_run_k_9);
	assign w_sys_tmp2367 = 32'sh00001b56;
	assign w_sys_tmp2371 = (w_sys_tmp2372 + r_run_k_9);
	assign w_sys_tmp2372 = 32'sh00001b76;
	assign w_sys_tmp2376 = (w_sys_tmp2377 + r_run_k_9);
	assign w_sys_tmp2377 = 32'sh00001bb7;
	assign w_sys_tmp2381 = (w_sys_tmp2382 + r_run_k_9);
	assign w_sys_tmp2382 = 32'sh00001bd7;
	assign w_sys_tmp2386 = (w_sys_tmp2387 + r_run_k_9);
	assign w_sys_tmp2387 = 32'sh00001bf7;
	assign w_sys_tmp2391 = (w_sys_tmp2392 + r_run_k_9);
	assign w_sys_tmp2392 = 32'sh00001c38;
	assign w_sys_tmp2396 = (w_sys_tmp2397 + r_run_k_9);
	assign w_sys_tmp2397 = 32'sh00001c58;
	assign w_sys_tmp2401 = (w_sys_tmp2402 + r_run_k_9);
	assign w_sys_tmp2402 = 32'sh00001c78;
	assign w_sys_tmp2406 = (w_sys_tmp2407 + r_run_k_9);
	assign w_sys_tmp2407 = 32'sh00001cb9;
	assign w_sys_tmp2411 = (w_sys_tmp2412 + r_run_k_9);
	assign w_sys_tmp2412 = 32'sh00001cd9;
	assign w_sys_tmp2416 = (w_sys_tmp2417 + r_run_k_9);
	assign w_sys_tmp2417 = 32'sh00001cf9;
	assign w_sys_tmp2421 = (w_sys_tmp2422 + r_run_k_9);
	assign w_sys_tmp2422 = 32'sh00001d3a;
	assign w_sys_tmp2426 = (w_sys_tmp2427 + r_run_k_9);
	assign w_sys_tmp2427 = 32'sh00001d5a;
	assign w_sys_tmp2431 = (w_sys_tmp2432 + r_run_k_9);
	assign w_sys_tmp2432 = 32'sh00001d7a;
	assign w_sys_tmp2436 = (w_sys_tmp2437 + r_run_k_9);
	assign w_sys_tmp2437 = 32'sh00001dbb;
	assign w_sys_tmp2441 = (w_sys_tmp2442 + r_run_k_9);
	assign w_sys_tmp2442 = 32'sh00001ddb;
	assign w_sys_tmp2446 = (w_sys_tmp2447 + r_run_k_9);
	assign w_sys_tmp2447 = 32'sh00001dfb;
	assign w_sys_tmp2451 = (w_sys_tmp2452 + r_run_k_9);
	assign w_sys_tmp2452 = 32'sh00001e3c;
	assign w_sys_tmp2456 = (w_sys_tmp2457 + r_run_k_9);
	assign w_sys_tmp2457 = 32'sh00001e5c;
	assign w_sys_tmp2461 = (w_sys_tmp2462 + r_run_k_9);
	assign w_sys_tmp2462 = 32'sh00001e7c;
	assign w_sys_tmp2466 = (w_sys_tmp2467 + r_run_k_9);
	assign w_sys_tmp2467 = 32'sh00001ebd;
	assign w_sys_tmp2471 = (w_sys_tmp2472 + r_run_k_9);
	assign w_sys_tmp2472 = 32'sh00001edd;
	assign w_sys_tmp2476 = (w_sys_tmp2477 + r_run_k_9);
	assign w_sys_tmp2477 = 32'sh00001efd;
	assign w_sys_tmp2481 = (w_sys_tmp2482 + r_run_k_9);
	assign w_sys_tmp2482 = 32'sh00001f3e;
	assign w_sys_tmp2486 = (w_sys_tmp2487 + r_run_k_9);
	assign w_sys_tmp2487 = 32'sh00001f5e;
	assign w_sys_tmp2491 = (w_sys_tmp2492 + r_run_k_9);
	assign w_sys_tmp2492 = 32'sh00001f7e;
	assign w_sys_tmp2496 = (w_sys_tmp2497 + r_run_k_9);
	assign w_sys_tmp2497 = 32'sh00001fbf;
	assign w_sys_tmp2501 = (w_sys_tmp2502 + r_run_k_9);
	assign w_sys_tmp2502 = 32'sh00001fdf;
	assign w_sys_tmp2506 = (w_sys_tmp2507 + r_run_k_9);
	assign w_sys_tmp2507 = 32'sh00001fff;
	assign w_sys_tmp2511 = (w_sys_tmp2512 + r_run_k_9);
	assign w_sys_tmp2512 = 32'sh00002040;
	assign w_sys_tmp2516 = (w_sys_tmp2517 + r_run_k_9);
	assign w_sys_tmp2517 = 32'sh00002060;
	assign w_sys_tmp2521 = (w_sys_tmp2522 + r_run_k_9);
	assign w_sys_tmp2522 = 32'sh00002080;
	assign w_sys_tmp2525 = (r_run_k_9 + w_sys_intOne);
	assign w_sys_tmp2526 = 32'sh00000041;
	assign w_sys_tmp2527 = ( !w_sys_tmp2528 );
	assign w_sys_tmp2528 = (w_sys_tmp2529 < r_run_k_9);
	assign w_sys_tmp2529 = 32'sh00000080;
	assign w_sys_tmp2532 = (w_sys_tmp2533 + r_run_k_9);
	assign w_sys_tmp2533 = 32'sh00000102;
	assign w_sys_tmp2534 = w_sub04_result_dataout;
	assign w_sys_tmp2538 = (w_sys_tmp2539 + r_run_k_9);
	assign w_sys_tmp2539 = 32'sh00000183;
	assign w_sys_tmp2544 = (w_sys_tmp2545 + r_run_k_9);
	assign w_sys_tmp2545 = 32'sh00000204;
	assign w_sys_tmp2550 = (w_sys_tmp2551 + r_run_k_9);
	assign w_sys_tmp2551 = 32'sh00000285;
	assign w_sys_tmp2556 = (w_sys_tmp2557 + r_run_k_9);
	assign w_sys_tmp2557 = 32'sh00000306;
	assign w_sys_tmp2562 = (w_sys_tmp2563 + r_run_k_9);
	assign w_sys_tmp2563 = 32'sh00000387;
	assign w_sys_tmp2568 = (w_sys_tmp2569 + r_run_k_9);
	assign w_sys_tmp2569 = 32'sh00000408;
	assign w_sys_tmp2574 = (w_sys_tmp2575 + r_run_k_9);
	assign w_sys_tmp2575 = 32'sh00000489;
	assign w_sys_tmp2580 = (w_sys_tmp2581 + r_run_k_9);
	assign w_sys_tmp2581 = 32'sh0000050a;
	assign w_sys_tmp2586 = (w_sys_tmp2587 + r_run_k_9);
	assign w_sys_tmp2587 = 32'sh0000058b;
	assign w_sys_tmp2592 = (w_sys_tmp2593 + r_run_k_9);
	assign w_sys_tmp2593 = 32'sh0000060c;
	assign w_sys_tmp2598 = (w_sys_tmp2599 + r_run_k_9);
	assign w_sys_tmp2599 = 32'sh0000068d;
	assign w_sys_tmp2604 = (w_sys_tmp2605 + r_run_k_9);
	assign w_sys_tmp2605 = 32'sh0000070e;
	assign w_sys_tmp2610 = (w_sys_tmp2611 + r_run_k_9);
	assign w_sys_tmp2611 = 32'sh0000078f;
	assign w_sys_tmp2616 = (w_sys_tmp2617 + r_run_k_9);
	assign w_sys_tmp2617 = 32'sh00000810;
	assign w_sys_tmp2622 = (w_sys_tmp2623 + r_run_k_9);
	assign w_sys_tmp2623 = 32'sh00000891;
	assign w_sys_tmp2628 = (w_sys_tmp2629 + r_run_k_9);
	assign w_sys_tmp2629 = 32'sh00000912;
	assign w_sys_tmp2634 = (w_sys_tmp2635 + r_run_k_9);
	assign w_sys_tmp2635 = 32'sh00000993;
	assign w_sys_tmp2640 = (w_sys_tmp2641 + r_run_k_9);
	assign w_sys_tmp2641 = 32'sh00000a14;
	assign w_sys_tmp2646 = (w_sys_tmp2647 + r_run_k_9);
	assign w_sys_tmp2647 = 32'sh00000a95;
	assign w_sys_tmp2652 = (w_sys_tmp2653 + r_run_k_9);
	assign w_sys_tmp2653 = 32'sh00000b16;
	assign w_sys_tmp2658 = (w_sys_tmp2659 + r_run_k_9);
	assign w_sys_tmp2659 = 32'sh00000b97;
	assign w_sys_tmp2664 = (w_sys_tmp2665 + r_run_k_9);
	assign w_sys_tmp2665 = 32'sh00000c18;
	assign w_sys_tmp2670 = (w_sys_tmp2671 + r_run_k_9);
	assign w_sys_tmp2671 = 32'sh00000c99;
	assign w_sys_tmp2676 = (w_sys_tmp2677 + r_run_k_9);
	assign w_sys_tmp2677 = 32'sh00000d1a;
	assign w_sys_tmp2682 = (w_sys_tmp2683 + r_run_k_9);
	assign w_sys_tmp2683 = 32'sh00000d9b;
	assign w_sys_tmp2688 = (w_sys_tmp2689 + r_run_k_9);
	assign w_sys_tmp2689 = 32'sh00000e1c;
	assign w_sys_tmp2694 = (w_sys_tmp2695 + r_run_k_9);
	assign w_sys_tmp2695 = 32'sh00000e9d;
	assign w_sys_tmp2700 = (w_sys_tmp2701 + r_run_k_9);
	assign w_sys_tmp2701 = 32'sh00000f1e;
	assign w_sys_tmp2706 = (w_sys_tmp2707 + r_run_k_9);
	assign w_sys_tmp2707 = 32'sh00000f9f;
	assign w_sys_tmp2712 = (w_sys_tmp2713 + r_run_k_9);
	assign w_sys_tmp2713 = 32'sh00001020;
	assign w_sys_tmp2718 = (w_sys_tmp2719 + r_run_k_9);
	assign w_sys_tmp2719 = 32'sh000010a1;
	assign w_sys_tmp2723 = (w_sys_tmp2724 + r_run_k_9);
	assign w_sys_tmp2724 = 32'sh000010c1;
	assign w_sys_tmp2728 = (w_sys_tmp2729 + r_run_k_9);
	assign w_sys_tmp2729 = 32'sh000010e1;
	assign w_sys_tmp2733 = (w_sys_tmp2734 + r_run_k_9);
	assign w_sys_tmp2734 = 32'sh00001122;
	assign w_sys_tmp2738 = (w_sys_tmp2739 + r_run_k_9);
	assign w_sys_tmp2739 = 32'sh00001142;
	assign w_sys_tmp2743 = (w_sys_tmp2744 + r_run_k_9);
	assign w_sys_tmp2744 = 32'sh00001162;
	assign w_sys_tmp2748 = (w_sys_tmp2749 + r_run_k_9);
	assign w_sys_tmp2749 = 32'sh000011a3;
	assign w_sys_tmp2753 = (w_sys_tmp2754 + r_run_k_9);
	assign w_sys_tmp2754 = 32'sh000011c3;
	assign w_sys_tmp2758 = (w_sys_tmp2759 + r_run_k_9);
	assign w_sys_tmp2759 = 32'sh000011e3;
	assign w_sys_tmp2763 = (w_sys_tmp2764 + r_run_k_9);
	assign w_sys_tmp2764 = 32'sh00001224;
	assign w_sys_tmp2768 = (w_sys_tmp2769 + r_run_k_9);
	assign w_sys_tmp2769 = 32'sh00001244;
	assign w_sys_tmp2773 = (w_sys_tmp2774 + r_run_k_9);
	assign w_sys_tmp2774 = 32'sh00001264;
	assign w_sys_tmp2778 = (w_sys_tmp2779 + r_run_k_9);
	assign w_sys_tmp2779 = 32'sh000012a5;
	assign w_sys_tmp2783 = (w_sys_tmp2784 + r_run_k_9);
	assign w_sys_tmp2784 = 32'sh000012c5;
	assign w_sys_tmp2788 = (w_sys_tmp2789 + r_run_k_9);
	assign w_sys_tmp2789 = 32'sh000012e5;
	assign w_sys_tmp2793 = (w_sys_tmp2794 + r_run_k_9);
	assign w_sys_tmp2794 = 32'sh00001326;
	assign w_sys_tmp2798 = (w_sys_tmp2799 + r_run_k_9);
	assign w_sys_tmp2799 = 32'sh00001346;
	assign w_sys_tmp2803 = (w_sys_tmp2804 + r_run_k_9);
	assign w_sys_tmp2804 = 32'sh00001366;
	assign w_sys_tmp2808 = (w_sys_tmp2809 + r_run_k_9);
	assign w_sys_tmp2809 = 32'sh000013a7;
	assign w_sys_tmp2813 = (w_sys_tmp2814 + r_run_k_9);
	assign w_sys_tmp2814 = 32'sh000013c7;
	assign w_sys_tmp2818 = (w_sys_tmp2819 + r_run_k_9);
	assign w_sys_tmp2819 = 32'sh000013e7;
	assign w_sys_tmp2823 = (w_sys_tmp2824 + r_run_k_9);
	assign w_sys_tmp2824 = 32'sh00001428;
	assign w_sys_tmp2828 = (w_sys_tmp2829 + r_run_k_9);
	assign w_sys_tmp2829 = 32'sh00001448;
	assign w_sys_tmp2833 = (w_sys_tmp2834 + r_run_k_9);
	assign w_sys_tmp2834 = 32'sh00001468;
	assign w_sys_tmp2838 = (w_sys_tmp2839 + r_run_k_9);
	assign w_sys_tmp2839 = 32'sh000014a9;
	assign w_sys_tmp2843 = (w_sys_tmp2844 + r_run_k_9);
	assign w_sys_tmp2844 = 32'sh000014c9;
	assign w_sys_tmp2848 = (w_sys_tmp2849 + r_run_k_9);
	assign w_sys_tmp2849 = 32'sh000014e9;
	assign w_sys_tmp2853 = (w_sys_tmp2854 + r_run_k_9);
	assign w_sys_tmp2854 = 32'sh0000152a;
	assign w_sys_tmp2858 = (w_sys_tmp2859 + r_run_k_9);
	assign w_sys_tmp2859 = 32'sh0000154a;
	assign w_sys_tmp2863 = (w_sys_tmp2864 + r_run_k_9);
	assign w_sys_tmp2864 = 32'sh0000156a;
	assign w_sys_tmp2868 = (w_sys_tmp2869 + r_run_k_9);
	assign w_sys_tmp2869 = 32'sh000015ab;
	assign w_sys_tmp2873 = (w_sys_tmp2874 + r_run_k_9);
	assign w_sys_tmp2874 = 32'sh000015cb;
	assign w_sys_tmp2878 = (w_sys_tmp2879 + r_run_k_9);
	assign w_sys_tmp2879 = 32'sh000015eb;
	assign w_sys_tmp2883 = (w_sys_tmp2884 + r_run_k_9);
	assign w_sys_tmp2884 = 32'sh0000162c;
	assign w_sys_tmp2888 = (w_sys_tmp2889 + r_run_k_9);
	assign w_sys_tmp2889 = 32'sh0000164c;
	assign w_sys_tmp2893 = (w_sys_tmp2894 + r_run_k_9);
	assign w_sys_tmp2894 = 32'sh0000166c;
	assign w_sys_tmp2898 = (w_sys_tmp2899 + r_run_k_9);
	assign w_sys_tmp2899 = 32'sh000016ad;
	assign w_sys_tmp2903 = (w_sys_tmp2904 + r_run_k_9);
	assign w_sys_tmp2904 = 32'sh000016cd;
	assign w_sys_tmp2908 = (w_sys_tmp2909 + r_run_k_9);
	assign w_sys_tmp2909 = 32'sh000016ed;
	assign w_sys_tmp2913 = (w_sys_tmp2914 + r_run_k_9);
	assign w_sys_tmp2914 = 32'sh0000172e;
	assign w_sys_tmp2918 = (w_sys_tmp2919 + r_run_k_9);
	assign w_sys_tmp2919 = 32'sh0000174e;
	assign w_sys_tmp2923 = (w_sys_tmp2924 + r_run_k_9);
	assign w_sys_tmp2924 = 32'sh0000176e;
	assign w_sys_tmp2928 = (w_sys_tmp2929 + r_run_k_9);
	assign w_sys_tmp2929 = 32'sh000017af;
	assign w_sys_tmp2933 = (w_sys_tmp2934 + r_run_k_9);
	assign w_sys_tmp2934 = 32'sh000017cf;
	assign w_sys_tmp2938 = (w_sys_tmp2939 + r_run_k_9);
	assign w_sys_tmp2939 = 32'sh000017ef;
	assign w_sys_tmp2943 = (w_sys_tmp2944 + r_run_k_9);
	assign w_sys_tmp2944 = 32'sh00001830;
	assign w_sys_tmp2948 = (w_sys_tmp2949 + r_run_k_9);
	assign w_sys_tmp2949 = 32'sh00001850;
	assign w_sys_tmp2953 = (w_sys_tmp2954 + r_run_k_9);
	assign w_sys_tmp2954 = 32'sh00001870;
	assign w_sys_tmp2958 = (w_sys_tmp2959 + r_run_k_9);
	assign w_sys_tmp2959 = 32'sh000018b1;
	assign w_sys_tmp2963 = (w_sys_tmp2964 + r_run_k_9);
	assign w_sys_tmp2964 = 32'sh000018d1;
	assign w_sys_tmp2968 = (w_sys_tmp2969 + r_run_k_9);
	assign w_sys_tmp2969 = 32'sh000018f1;
	assign w_sys_tmp2973 = (w_sys_tmp2974 + r_run_k_9);
	assign w_sys_tmp2974 = 32'sh00001932;
	assign w_sys_tmp2978 = (w_sys_tmp2979 + r_run_k_9);
	assign w_sys_tmp2979 = 32'sh00001952;
	assign w_sys_tmp2983 = (w_sys_tmp2984 + r_run_k_9);
	assign w_sys_tmp2984 = 32'sh00001972;
	assign w_sys_tmp2988 = (w_sys_tmp2989 + r_run_k_9);
	assign w_sys_tmp2989 = 32'sh000019b3;
	assign w_sys_tmp2993 = (w_sys_tmp2994 + r_run_k_9);
	assign w_sys_tmp2994 = 32'sh000019d3;
	assign w_sys_tmp2998 = (w_sys_tmp2999 + r_run_k_9);
	assign w_sys_tmp2999 = 32'sh000019f3;
	assign w_sys_tmp3003 = (w_sys_tmp3004 + r_run_k_9);
	assign w_sys_tmp3004 = 32'sh00001a34;
	assign w_sys_tmp3008 = (w_sys_tmp3009 + r_run_k_9);
	assign w_sys_tmp3009 = 32'sh00001a54;
	assign w_sys_tmp3013 = (w_sys_tmp3014 + r_run_k_9);
	assign w_sys_tmp3014 = 32'sh00001a74;
	assign w_sys_tmp3018 = (w_sys_tmp3019 + r_run_k_9);
	assign w_sys_tmp3019 = 32'sh00001ab5;
	assign w_sys_tmp3023 = (w_sys_tmp3024 + r_run_k_9);
	assign w_sys_tmp3024 = 32'sh00001ad5;
	assign w_sys_tmp3028 = (w_sys_tmp3029 + r_run_k_9);
	assign w_sys_tmp3029 = 32'sh00001af5;
	assign w_sys_tmp3033 = (w_sys_tmp3034 + r_run_k_9);
	assign w_sys_tmp3034 = 32'sh00001b36;
	assign w_sys_tmp3038 = (w_sys_tmp3039 + r_run_k_9);
	assign w_sys_tmp3039 = 32'sh00001b56;
	assign w_sys_tmp3043 = (w_sys_tmp3044 + r_run_k_9);
	assign w_sys_tmp3044 = 32'sh00001b76;
	assign w_sys_tmp3048 = (w_sys_tmp3049 + r_run_k_9);
	assign w_sys_tmp3049 = 32'sh00001bb7;
	assign w_sys_tmp3053 = (w_sys_tmp3054 + r_run_k_9);
	assign w_sys_tmp3054 = 32'sh00001bd7;
	assign w_sys_tmp3058 = (w_sys_tmp3059 + r_run_k_9);
	assign w_sys_tmp3059 = 32'sh00001bf7;
	assign w_sys_tmp3063 = (w_sys_tmp3064 + r_run_k_9);
	assign w_sys_tmp3064 = 32'sh00001c38;
	assign w_sys_tmp3068 = (w_sys_tmp3069 + r_run_k_9);
	assign w_sys_tmp3069 = 32'sh00001c58;
	assign w_sys_tmp3073 = (w_sys_tmp3074 + r_run_k_9);
	assign w_sys_tmp3074 = 32'sh00001c78;
	assign w_sys_tmp3078 = (w_sys_tmp3079 + r_run_k_9);
	assign w_sys_tmp3079 = 32'sh00001cb9;
	assign w_sys_tmp3083 = (w_sys_tmp3084 + r_run_k_9);
	assign w_sys_tmp3084 = 32'sh00001cd9;
	assign w_sys_tmp3088 = (w_sys_tmp3089 + r_run_k_9);
	assign w_sys_tmp3089 = 32'sh00001cf9;
	assign w_sys_tmp3093 = (w_sys_tmp3094 + r_run_k_9);
	assign w_sys_tmp3094 = 32'sh00001d3a;
	assign w_sys_tmp3098 = (w_sys_tmp3099 + r_run_k_9);
	assign w_sys_tmp3099 = 32'sh00001d5a;
	assign w_sys_tmp3103 = (w_sys_tmp3104 + r_run_k_9);
	assign w_sys_tmp3104 = 32'sh00001d7a;
	assign w_sys_tmp3108 = (w_sys_tmp3109 + r_run_k_9);
	assign w_sys_tmp3109 = 32'sh00001dbb;
	assign w_sys_tmp3113 = (w_sys_tmp3114 + r_run_k_9);
	assign w_sys_tmp3114 = 32'sh00001ddb;
	assign w_sys_tmp3118 = (w_sys_tmp3119 + r_run_k_9);
	assign w_sys_tmp3119 = 32'sh00001dfb;
	assign w_sys_tmp3123 = (w_sys_tmp3124 + r_run_k_9);
	assign w_sys_tmp3124 = 32'sh00001e3c;
	assign w_sys_tmp3128 = (w_sys_tmp3129 + r_run_k_9);
	assign w_sys_tmp3129 = 32'sh00001e5c;
	assign w_sys_tmp3133 = (w_sys_tmp3134 + r_run_k_9);
	assign w_sys_tmp3134 = 32'sh00001e7c;
	assign w_sys_tmp3138 = (w_sys_tmp3139 + r_run_k_9);
	assign w_sys_tmp3139 = 32'sh00001ebd;
	assign w_sys_tmp3143 = (w_sys_tmp3144 + r_run_k_9);
	assign w_sys_tmp3144 = 32'sh00001edd;
	assign w_sys_tmp3148 = (w_sys_tmp3149 + r_run_k_9);
	assign w_sys_tmp3149 = 32'sh00001efd;
	assign w_sys_tmp3153 = (w_sys_tmp3154 + r_run_k_9);
	assign w_sys_tmp3154 = 32'sh00001f3e;
	assign w_sys_tmp3158 = (w_sys_tmp3159 + r_run_k_9);
	assign w_sys_tmp3159 = 32'sh00001f5e;
	assign w_sys_tmp3163 = (w_sys_tmp3164 + r_run_k_9);
	assign w_sys_tmp3164 = 32'sh00001f7e;
	assign w_sys_tmp3168 = (w_sys_tmp3169 + r_run_k_9);
	assign w_sys_tmp3169 = 32'sh00001fbf;
	assign w_sys_tmp3173 = (w_sys_tmp3174 + r_run_k_9);
	assign w_sys_tmp3174 = 32'sh00001fdf;
	assign w_sys_tmp3178 = (w_sys_tmp3179 + r_run_k_9);
	assign w_sys_tmp3179 = 32'sh00001fff;
	assign w_sys_tmp3183 = (w_sys_tmp3184 + r_run_k_9);
	assign w_sys_tmp3184 = 32'sh00002040;
	assign w_sys_tmp3188 = (w_sys_tmp3189 + r_run_k_9);
	assign w_sys_tmp3189 = 32'sh00002060;
	assign w_sys_tmp3193 = (w_sys_tmp3194 + r_run_k_9);
	assign w_sys_tmp3194 = 32'sh00002080;
	assign w_sys_tmp3197 = (r_run_k_9 + w_sys_intOne);
	assign w_sys_tmp3198 = w_fld_u_0_dataout_1;
	assign w_sys_tmp3199 = 32'sh000000dc;


	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_result_1_addr_0 (w_sub05_result_addr),
			.i_fld_result_1_datain_0 (w_sub05_result_datain),
			.o_fld_result_1_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h37: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_return <= 32'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h34: begin
							r_sys_run_return <= r_sys_tmp0_float;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_phase <= 6'h2;
						end

						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h4;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8) ? 6'h9 : 6'hf);

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h5;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11) ? 6'hd : 6'h6);

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_run_phase <= 6'ha;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp56) ? 6'h14 : 6'h35);

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h10;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp59) ? 6'h18 : 6'h1a);

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sys_run_phase <= 6'h15;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp223) ? 6'h1e : 6'h20);

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h88)) begin
										r_sys_run_phase <= 6'h1b;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1039) ? 6'h24 : 6'h25);

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h88)) begin
										r_sys_run_phase <= 6'h21;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_phase <= 6'h27;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								4'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_phase <= 6'h29;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1855) ? 6'h2d : 6'h2f);

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h80)) begin
										r_sys_run_phase <= 6'h2a;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2527) ? 6'h33 : 6'h11);

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h80)) begin
										r_sys_run_phase <= 6'h30;

									end
								end

							endcase
						end

						6'h34: begin
							r_sys_run_phase <= 6'h37;
						end

						6'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_run_phase <= 6'h34;

									end
								end

							endcase
						end

						6'h37: begin
							r_sys_run_phase <= 6'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h88)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h88)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h80)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h80)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						6'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 8'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h88)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h87)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h88)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h87)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						6'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h7f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h7f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

						6'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h1)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sys_run_step <= 8'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						6'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						6'h37: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp15[14:0] );

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp77[14:0] );

									end
									else
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp67[14:0] );

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp63[14:0] );

									end
									else
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp72[14:0] );

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h77)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp942[14:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp900[14:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp654[14:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp540[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp378[14:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp642[14:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp660[14:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp522[14:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp762[14:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp840[14:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp564[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp324[14:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp684[14:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp510[14:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp534[14:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp786[14:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp636[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp270[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp408[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp306[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp342[14:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp756[14:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp948[14:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp798[14:0] );

									end
									else
									if((r_sys_run_step==8'h20) || (r_sys_run_step==8'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp420[14:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp702[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp330[14:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp486[14:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp678[14:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp882[14:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp774[14:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp750[14:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp606[14:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp570[14:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp984[14:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp816[14:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp834[14:0] );

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1032[14:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp558[14:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp894[14:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp516[14:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp858[14:0] );

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp972[14:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp588[14:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp936[14:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp480[14:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp708[14:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp234[14:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp888[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp318[14:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp672[14:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp648[14:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp852[14:0] );

									end
									else
									if((r_sys_run_step==8'h85)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1026[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp384[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp372[14:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp462[14:0] );

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1014[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp258[14:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp846[14:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp492[14:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp924[14:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp450[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp294[14:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1008[14:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp690[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp240[14:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp714[14:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp732[14:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp930[14:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp906[14:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp768[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp336[14:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp744[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp288[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp360[14:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp546[14:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp696[14:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp228[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp414[14:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp864[14:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp456[14:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp720[14:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp576[14:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp804[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp276[14:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp870[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp402[14:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp498[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp300[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp264[14:0] );

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp978[14:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp918[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp282[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp354[14:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp474[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp252[14:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp780[14:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1002[14:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp438[14:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp612[14:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp468[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp390[14:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp600[14:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp552[14:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp876[14:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp432[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp246[14:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp990[14:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp810[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp396[14:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp792[14:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp912[14:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp528[14:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp630[14:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp954[14:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp822[14:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp966[14:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp594[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp348[14:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp504[14:0] );

									end
									else
									if((r_sys_run_step==8'h84)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1020[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp312[14:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp582[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp366[14:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp618[14:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp996[14:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp666[14:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp726[14:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp738[14:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp960[14:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp828[14:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp624[14:0] );

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1188[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1140[14:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1596[14:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1338[14:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1446[14:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1440[14:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1332[14:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1572[14:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1602[14:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1290[14:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1686[14:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1764[14:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1728[14:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1680[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1194[14:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1482[14:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1626[14:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1800[14:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1452[14:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1590[14:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1368[14:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1734[14:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1296[14:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1272[14:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1464[14:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1374[14:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1776[14:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1656[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1098[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1092[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1062[14:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1566[14:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1638[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1056[14:0] );

									end
									else
									if((r_sys_run_step==8'h85)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1842[14:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1050[14:0] );

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1848[14:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1644[14:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1632[14:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1512[14:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1524[14:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1698[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1164[14:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1584[14:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1458[14:0] );

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1794[14:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1746[14:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1488[14:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1362[14:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1740[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1182[14:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1620[14:0] );

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1788[14:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1494[14:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1668[14:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1356[14:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1320[14:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1530[14:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1818[14:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1254[14:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1812[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1212[14:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1770[14:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1278[14:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1542[14:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1044[14:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1470[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1086[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1110[14:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1710[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1068[14:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1560[14:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1302[14:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1428[14:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1326[14:0] );

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1830[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1218[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1116[14:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1434[14:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1548[14:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1248[14:0] );

									end
									else
									if((r_sys_run_step==8'h20) || (r_sys_run_step==8'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1236[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1200[14:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1722[14:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1758[14:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1266[14:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1422[14:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1782[14:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1404[14:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1476[14:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1518[14:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1614[14:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1350[14:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1806[14:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1692[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1074[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1128[14:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1824[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1170[14:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1536[14:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1500[14:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1608[14:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1308[14:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1578[14:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1380[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1176[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1134[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1122[14:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1674[14:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1662[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f) || (r_sys_run_step==8'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1230[14:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1704[14:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1392[14:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1554[14:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1752[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1158[14:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1410[14:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1716[14:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1344[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1146[14:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1386[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1206[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1152[14:0] );

									end
									else
									if((r_sys_run_step==8'h84)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1836[14:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1284[14:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1314[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1224[14:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1506[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1080[14:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1398[14:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1416[14:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1650[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1104[14:0] );

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1896[14:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2316[14:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2426[14:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2346[14:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2476[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2004[14:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2286[14:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2051[14:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2251[14:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2496[14:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2381[14:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2081[14:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2141[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2034[14:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2296[14:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2361[14:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2121[14:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2371[14:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2091[14:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2511[14:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2086[14:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2061[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1866[14:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2416[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2016[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1926[14:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2246[14:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2111[14:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2291[14:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2226[14:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2231[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1980[14:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2321[14:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2336[14:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2171[14:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2146[14:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2446[14:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2241[14:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2266[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1992[14:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2151[14:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2186[14:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2256[14:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2516[14:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2521[14:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2401[14:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2421[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1872[14:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2441[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2022[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2028[14:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2456[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1890[14:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2351[14:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2106[14:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2466[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1962[14:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2461[14:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2326[14:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2391[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2010[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1950[14:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2276[14:0] );

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2501[14:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2301[14:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2196[14:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2436[14:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2261[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1944[14:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2191[14:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2166[14:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2481[14:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2271[14:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2071[14:0] );

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2506[14:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2131[14:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2101[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1884[14:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2201[14:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2341[14:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2491[14:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2376[14:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2136[14:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2211[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1878[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1908[14:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2281[14:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2366[14:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2451[14:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2046[14:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2161[14:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2306[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1914[14:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2221[14:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2331[14:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2406[14:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2096[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1932[14:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2431[14:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2486[14:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2040[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1974[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1968[14:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2311[14:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2076[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1902[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1998[14:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2126[14:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2386[14:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2176[14:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2156[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1956[14:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2181[14:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2216[14:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2471[14:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2411[14:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2206[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1920[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1860[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1938[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1986[14:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2396[14:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2056[14:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2236[14:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2066[14:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2356[14:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2116[14:0] );

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h43)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2888[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2586[14:0] );

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3178[14:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3098[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2682[14:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3083[14:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2898[14:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3063[14:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2853[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2610[14:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2983[14:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3023[14:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2903[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2694[14:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3043[14:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2833[14:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2883[14:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2848[14:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2878[14:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3058[14:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3048[14:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3093[14:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2803[14:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3113[14:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2828[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2592[14:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2723[14:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2813[14:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3053[14:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2908[14:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2933[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2604[14:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2958[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2658[14:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3183[14:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3118[14:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3003[14:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2712[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2700[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2688[14:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2943[14:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3143[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2574[14:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2948[14:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2913[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2568[14:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3123[14:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2763[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2652[14:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3033[14:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3163[14:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3138[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2532[14:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2918[14:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2793[14:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3193[14:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2768[14:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2968[14:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2928[14:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2858[14:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2728[14:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3148[14:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2863[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2544[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2664[14:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3188[14:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2778[14:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2753[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2556[14:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3028[14:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2718[14:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3038[14:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2823[14:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2868[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2646[14:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3133[14:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2773[14:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2808[14:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3168[14:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3013[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2538[14:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3158[14:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2748[14:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2973[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2616[14:0] );

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3173[14:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2798[14:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2873[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2640[14:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3103[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2634[14:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2953[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2622[14:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2743[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2706[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2562[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2676[14:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2963[14:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2993[14:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2988[14:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3153[14:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2978[14:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2838[14:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3108[14:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3068[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2670[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2598[14:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2843[14:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3128[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2550[14:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2738[14:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2733[14:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2938[14:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2998[14:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3073[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2628[14:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2818[14:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2893[14:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3078[14:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2783[14:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2923[14:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3088[14:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3008[14:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2788[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2580[14:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3018[14:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2758[14:0] );

									end
								end

							endcase
						end

						6'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp3199[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1a)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp75;

									end
									else
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h3) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h19) || (r_sys_run_step==8'h1b)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp70;

									end
									else
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h18)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp65;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h5a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp82_float;

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp76_float;

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp74_float;

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h20)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp1862;

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp77_float;

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp87_float;

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp81_float;

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp90_float;

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp85_float;

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp91_float;

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp83_float;

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp92_float;

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp75_float;

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp93_float;

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp84_float;

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp89_float;

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp80_float;

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp88_float;

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp78_float;

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==8'h21) || (r_sys_run_step==8'h7e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp94_float;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h5e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp82_float;

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h20)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp2534;

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp76_float;

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp74_float;

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp77_float;

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp87_float;

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp81_float;

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp90_float;

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp85_float;

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp91_float;

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp83_float;

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp92_float;

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp75_float;

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp93_float;

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp84_float;

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp89_float;

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp80_float;

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp88_float;

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp78_float;

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==8'h21) || (r_sys_run_step==8'h7e)) begin
										r_fld_u_0_datain_1 <= r_sys_tmp94_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1b)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h86)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h80)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h80)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_9 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_9 <= w_sys_tmp10;

									end
								end

							endcase
						end

						6'h1a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_9 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h88)) begin
										r_run_k_9 <= w_sys_tmp1037;

									end
								end

							endcase
						end

						6'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_9 <= w_sys_tmp1038;

									end
								end

							endcase
						end

						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h88)) begin
										r_run_k_9 <= w_sys_tmp1853;

									end
								end

							endcase
						end

						6'h29: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_9 <= w_sys_tmp1854;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h80)) begin
										r_run_k_9 <= w_sys_tmp2525;

									end
								end

							endcase
						end

						6'h2f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_k_9 <= w_sys_tmp2526;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h80)) begin
										r_run_k_9 <= w_sys_tmp3197;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_10 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h6)) begin
										r_run_j_10 <= w_sys_tmp19;

									end
								end

							endcase
						end

						6'h14: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_j_10 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0) || (r_sys_run_step==8'h4) || (r_sys_run_step==8'h8) || (r_sys_run_step==8'hc) || (r_sys_run_step==8'h10) || (r_sys_run_step==8'h14) || (r_sys_run_step==8'h18)) begin
										r_run_j_10 <= w_sys_tmp84;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_n_11 <= w_sys_intOne;

									end
								end

							endcase
						end

						6'h11: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_n_11 <= w_sys_tmp58;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_mx_12 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_my_13 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_nlast_14 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dx_15 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dy_16 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_dt_17 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r1_18 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_r2_19 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy0_j_20 <= r_run_j_10;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h3) || (r_sys_run_step==8'h7) || (r_sys_run_step==8'hb) || (r_sys_run_step==8'hf) || (r_sys_run_step==8'h13) || (r_sys_run_step==8'h17) || (r_sys_run_step==8'h1b)) begin
										r_run_copy0_j_20 <= w_sys_tmp81;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy1_j_21 <= r_run_j_10;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h6) || (r_sys_run_step==8'ha) || (r_sys_run_step==8'he) || (r_sys_run_step==8'h12) || (r_sys_run_step==8'h16) || (r_sys_run_step==8'h1a)) begin
										r_run_copy1_j_21 <= w_sys_tmp82;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h14: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_run_copy2_j_22 <= r_run_j_10;

									end
								end

							endcase
						end

						6'h18: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1) || (r_sys_run_step==8'h5) || (r_sys_run_step==8'h9) || (r_sys_run_step==8'hd) || (r_sys_run_step==8'h11) || (r_sys_run_step==8'h15) || (r_sys_run_step==8'h19)) begin
										r_run_copy2_j_22 <= w_sys_tmp83;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h88)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp1032[14:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp942[14:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp780[14:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp654[14:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp906[14:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp744[14:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp438[14:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp546[14:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp762[14:0] );

									end
									else
									if((r_sys_run_step==8'h3a)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp564[14:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp600[14:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp510[14:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp456[14:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp636[14:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp708[14:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp888[14:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp672[14:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp852[14:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp870[14:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp528[14:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp798[14:0] );

									end
									else
									if((r_sys_run_step==8'h85)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp1014[14:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp492[14:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp582[14:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp924[14:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp978[14:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp618[14:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp474[14:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp816[14:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp996[14:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp690[14:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp726[14:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp834[14:0] );

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp960[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h88)) begin
										r_sub03_u_datain <= w_sys_tmp230;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h88)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2461[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2326[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2281[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2161[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2476[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2221[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2431[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2146[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2446[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2251[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2266[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2311[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2191[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2386[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2176[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2521[14:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2071[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2401[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2296[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2506[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2131[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2206[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2371[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2086[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2101[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2341[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2416[14:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2056[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2236[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2491[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2356[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2116[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1f)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h39)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp558[14:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp900[14:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp540[14:0] );

									end
									else
									if((r_sys_run_step==8'h33)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp522[14:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp612[14:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp468[14:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp684[14:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp972[14:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp432[14:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp864[14:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp936[14:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp720[14:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp990[14:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp810[14:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp756[14:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp576[14:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp648[14:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp792[14:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp1026[14:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp702[14:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp630[14:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp954[14:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp486[14:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp882[14:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp594[14:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp774[14:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp846[14:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp504[14:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp918[14:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp450[14:0] );

									end
									else
									if((r_sys_run_step==8'h84)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp1008[14:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp666[14:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp738[14:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp828[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h87)) begin
										r_sub02_u_datain <= w_sys_tmp230;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h87)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2231[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2366[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2321[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2426[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2306[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2336[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2096[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2276[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2486[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2171[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2501[14:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2051[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2381[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2261[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2126[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2186[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2081[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2516[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2156[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2216[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2141[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2471[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2441[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2411[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2456[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2201[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2246[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2396[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2351[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2111[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2291[14:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2066[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1f)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h53)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp714[14:0] );

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp1002[14:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp894[14:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp732[14:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp930[14:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp768[14:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp642[14:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp660[14:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp516[14:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp840[14:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp858[14:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp696[14:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp552[14:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp534[14:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp414[14:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp876[14:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp588[14:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp786[14:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp480[14:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp804[14:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp948[14:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp912[14:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp498[14:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp420[14:0] );

									end
									else
									if((r_sys_run_step==8'h65)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp822[14:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp678[14:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp462[14:0] );

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp966[14:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp750[14:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp606[14:0] );

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp1020[14:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp570[14:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp984[14:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp624[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h23) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h86)) begin
										r_sub01_u_datain <= w_sys_tmp230;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h23) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h86)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hb)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2211[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2391[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2451[14:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2046[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2316[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2346[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2331[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2406[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2286[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2241[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2301[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2496[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2196[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2436[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2076[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2151[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2166[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2256[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2481[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2271[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2181[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2421[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2361[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2121[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2091[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2511[14:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2061[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2106[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2466[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2226[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2136[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2376[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1f)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp240[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp378[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp336[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp288[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp360[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp324[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp228[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp390[14:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp414[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp246[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp270[14:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp408[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp234[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp306[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp342[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp318[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp396[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp276[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp402[14:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp420[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp384[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp330[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp372[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp258[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp348[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp300[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp264[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp312[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp366[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp282[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp354[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp294[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp252[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h22)) begin
										r_sub00_u_datain <= w_sys_tmp230;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h1e: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h22)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1878[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1980[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1908[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1896[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2010[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1950[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1914[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1932[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2004[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2040[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1974[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1968[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1902[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1998[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1944[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1992[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1956[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2034[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1872[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1920[14:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1860[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1938[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2022[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1986[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1884[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2028[14:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1866[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2016[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1926[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1890[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp1962[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1e)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h3a)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1380[14:0] );

									end
									else
									if((r_sys_run_step==8'h55)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1542[14:0] );

									end
									else
									if((r_sys_run_step==8'h5e)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1596[14:0] );

									end
									else
									if((r_sys_run_step==8'h49)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1470[14:0] );

									end
									else
									if((r_sys_run_step==8'h88)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1848[14:0] );

									end
									else
									if((r_sys_run_step==8'h64)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1632[14:0] );

									end
									else
									if((r_sys_run_step==8'h2b)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1290[14:0] );

									end
									else
									if((r_sys_run_step==8'h52)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1524[14:0] );

									end
									else
									if((r_sys_run_step==8'h6d)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1686[14:0] );

									end
									else
									if((r_sys_run_step==8'h58)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1560[14:0] );

									end
									else
									if((r_sys_run_step==8'h70)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1704[14:0] );

									end
									else
									if((r_sys_run_step==8'h31)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1326[14:0] );

									end
									else
									if((r_sys_run_step==8'h85)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1830[14:0] );

									end
									else
									if((r_sys_run_step==8'h43)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1434[14:0] );

									end
									else
									if((r_sys_run_step==8'h7f)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1794[14:0] );

									end
									else
									if((r_sys_run_step==8'h4c)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1488[14:0] );

									end
									else
									if((r_sys_run_step==8'h46)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1452[14:0] );

									end
									else
									if((r_sys_run_step==8'h73)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1722[14:0] );

									end
									else
									if((r_sys_run_step==8'h34)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1344[14:0] );

									end
									else
									if((r_sys_run_step==8'h37)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1362[14:0] );

									end
									else
									if((r_sys_run_step==8'h76)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1740[14:0] );

									end
									else
									if((r_sys_run_step==8'h79)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1758[14:0] );

									end
									else
									if((r_sys_run_step==8'h28)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1272[14:0] );

									end
									else
									if((r_sys_run_step==8'h7c)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1776[14:0] );

									end
									else
									if((r_sys_run_step==8'h6a)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1668[14:0] );

									end
									else
									if((r_sys_run_step==8'h61)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1614[14:0] );

									end
									else
									if((r_sys_run_step==8'h25)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1254[14:0] );

									end
									else
									if((r_sys_run_step==8'h82)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1812[14:0] );

									end
									else
									if((r_sys_run_step==8'h4f)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1506[14:0] );

									end
									else
									if((r_sys_run_step==8'h40)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1416[14:0] );

									end
									else
									if((r_sys_run_step==8'h3d)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1398[14:0] );

									end
									else
									if((r_sys_run_step==8'h2e)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1308[14:0] );

									end
									else
									if((r_sys_run_step==8'h67)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1650[14:0] );

									end
									else
									if((r_sys_run_step==8'h5b)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp1578[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h88)) begin
										r_sub07_u_datain <= w_sys_tmp1046;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h25) || (r_sys_run_step==8'h28) || (r_sys_run_step==8'h2b) || (r_sys_run_step==8'h2e) || (r_sys_run_step==8'h31) || (r_sys_run_step==8'h34) || (r_sys_run_step==8'h37) || (r_sys_run_step==8'h3a) || (r_sys_run_step==8'h3d) || (r_sys_run_step==8'h40) || (r_sys_run_step==8'h43) || (r_sys_run_step==8'h46) || (r_sys_run_step==8'h49) || (r_sys_run_step==8'h4c) || (r_sys_run_step==8'h4f) || (r_sys_run_step==8'h52) || (r_sys_run_step==8'h55) || (r_sys_run_step==8'h58) || (r_sys_run_step==8'h5b) || (r_sys_run_step==8'h5e) || (r_sys_run_step==8'h61) || (r_sys_run_step==8'h64) || (r_sys_run_step==8'h67) || (r_sys_run_step==8'h6a) || (r_sys_run_step==8'h6d) || (r_sys_run_step==8'h70) || (r_sys_run_step==8'h73) || (r_sys_run_step==8'h76) || (r_sys_run_step==8'h79) || (r_sys_run_step==8'h7c) || (r_sys_run_step==8'h7f) || (r_sys_run_step==8'h82) || (r_sys_run_step==8'h85) || (r_sys_run_step==8'h88)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2908[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3178[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3118[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3028[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2983[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3133[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2773[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2938[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2833[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3043[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2998[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3073[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2893[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2818[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3013[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3163[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2848[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3193[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2923[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2878[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3058[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3103[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3088[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2788[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2953[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2968[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2803[14:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2743[14:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2728[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp3148[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2863[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2758[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1f)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h33)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1338[14:0] );

									end
									else
									if((r_sys_run_step==8'h45)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1446[14:0] );

									end
									else
									if((r_sys_run_step==8'h87)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1842[14:0] );

									end
									else
									if((r_sys_run_step==8'h66)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1644[14:0] );

									end
									else
									if((r_sys_run_step==8'h5a)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1572[14:0] );

									end
									else
									if((r_sys_run_step==8'h6f)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1698[14:0] );

									end
									else
									if((r_sys_run_step==8'h69)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1662[14:0] );

									end
									else
									if((r_sys_run_step==8'h42)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1428[14:0] );

									end
									else
									if((r_sys_run_step==8'h2d)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1302[14:0] );

									end
									else
									if((r_sys_run_step==8'h3c)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1392[14:0] );

									end
									else
									if((r_sys_run_step==8'h6c)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1680[14:0] );

									end
									else
									if((r_sys_run_step==8'h57)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1554[14:0] );

									end
									else
									if((r_sys_run_step==8'h78)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1752[14:0] );

									end
									else
									if((r_sys_run_step==8'h24)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1248[14:0] );

									end
									else
									if((r_sys_run_step==8'h4b)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1482[14:0] );

									end
									else
									if((r_sys_run_step==8'h63)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1626[14:0] );

									end
									else
									if((r_sys_run_step==8'h3f)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1410[14:0] );

									end
									else
									if((r_sys_run_step==8'h72)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1716[14:0] );

									end
									else
									if((r_sys_run_step==8'h5d)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1590[14:0] );

									end
									else
									if((r_sys_run_step==8'h75)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1734[14:0] );

									end
									else
									if((r_sys_run_step==8'h27)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1266[14:0] );

									end
									else
									if((r_sys_run_step==8'h48)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1464[14:0] );

									end
									else
									if((r_sys_run_step==8'h7e)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1788[14:0] );

									end
									else
									if((r_sys_run_step==8'h39)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1374[14:0] );

									end
									else
									if((r_sys_run_step==8'h36)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1356[14:0] );

									end
									else
									if((r_sys_run_step==8'h51)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1518[14:0] );

									end
									else
									if((r_sys_run_step==8'h30)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1320[14:0] );

									end
									else
									if((r_sys_run_step==8'h2a)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1284[14:0] );

									end
									else
									if((r_sys_run_step==8'h81)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1806[14:0] );

									end
									else
									if((r_sys_run_step==8'h7b)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1770[14:0] );

									end
									else
									if((r_sys_run_step==8'h84)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1824[14:0] );

									end
									else
									if((r_sys_run_step==8'h54)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1536[14:0] );

									end
									else
									if((r_sys_run_step==8'h4e)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1500[14:0] );

									end
									else
									if((r_sys_run_step==8'h60)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp1608[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h87)) begin
										r_sub06_u_datain <= w_sys_tmp1046;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h24) || (r_sys_run_step==8'h27) || (r_sys_run_step==8'h2a) || (r_sys_run_step==8'h2d) || (r_sys_run_step==8'h30) || (r_sys_run_step==8'h33) || (r_sys_run_step==8'h36) || (r_sys_run_step==8'h39) || (r_sys_run_step==8'h3c) || (r_sys_run_step==8'h3f) || (r_sys_run_step==8'h42) || (r_sys_run_step==8'h45) || (r_sys_run_step==8'h48) || (r_sys_run_step==8'h4b) || (r_sys_run_step==8'h4e) || (r_sys_run_step==8'h51) || (r_sys_run_step==8'h54) || (r_sys_run_step==8'h57) || (r_sys_run_step==8'h5a) || (r_sys_run_step==8'h5d) || (r_sys_run_step==8'h60) || (r_sys_run_step==8'h63) || (r_sys_run_step==8'h66) || (r_sys_run_step==8'h69) || (r_sys_run_step==8'h6c) || (r_sys_run_step==8'h6f) || (r_sys_run_step==8'h72) || (r_sys_run_step==8'h75) || (r_sys_run_step==8'h78) || (r_sys_run_step==8'h7b) || (r_sys_run_step==8'h7e) || (r_sys_run_step==8'h81) || (r_sys_run_step==8'h84) || (r_sys_run_step==8'h87)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2813[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3053[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2888[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2933[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3188[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2963[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3098[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2753[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2993[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2978[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3038[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3083[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3023[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3143[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3068[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2948[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2843[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3128[14:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2738[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2903[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2918[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3158[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2783[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3173[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2873[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2798[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2768[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3008[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2858[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp3113[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2828[14:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2723[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1f)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h65)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1638[14:0] );

									end
									else
									if((r_sys_run_step==8'h44)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1440[14:0] );

									end
									else
									if((r_sys_run_step==8'h32)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1332[14:0] );

									end
									else
									if((r_sys_run_step==8'h50)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1512[14:0] );

									end
									else
									if((r_sys_run_step==8'h5f)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1602[14:0] );

									end
									else
									if((r_sys_run_step==8'h71)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1710[14:0] );

									end
									else
									if((r_sys_run_step==8'h6b)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1674[14:0] );

									end
									else
									if((r_sys_run_step==8'h23)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1230[14:0] );

									end
									else
									if((r_sys_run_step==8'h7a)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1764[14:0] );

									end
									else
									if((r_sys_run_step==8'h5c)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1584[14:0] );

									end
									else
									if((r_sys_run_step==8'h74)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1728[14:0] );

									end
									else
									if((r_sys_run_step==8'h47)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1458[14:0] );

									end
									else
									if((r_sys_run_step==8'h56)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1548[14:0] );

									end
									else
									if((r_sys_run_step==8'h77)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1746[14:0] );

									end
									else
									if((r_sys_run_step==8'h80)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1800[14:0] );

									end
									else
									if((r_sys_run_step==8'h26)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1236[14:0] );

									end
									else
									if((r_sys_run_step==8'h3b)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1386[14:0] );

									end
									else
									if((r_sys_run_step==8'h38)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1368[14:0] );

									end
									else
									if((r_sys_run_step==8'h62)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1620[14:0] );

									end
									else
									if((r_sys_run_step==8'h2c)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1296[14:0] );

									end
									else
									if((r_sys_run_step==8'h41)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1422[14:0] );

									end
									else
									if((r_sys_run_step==8'h86)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1836[14:0] );

									end
									else
									if((r_sys_run_step==8'h7d)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1782[14:0] );

									end
									else
									if((r_sys_run_step==8'h4d)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1494[14:0] );

									end
									else
									if((r_sys_run_step==8'h3e)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1404[14:0] );

									end
									else
									if((r_sys_run_step==8'h4a)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1476[14:0] );

									end
									else
									if((r_sys_run_step==8'h68)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1656[14:0] );

									end
									else
									if((r_sys_run_step==8'h53)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1530[14:0] );

									end
									else
									if((r_sys_run_step==8'h83)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1818[14:0] );

									end
									else
									if((r_sys_run_step==8'h35)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1350[14:0] );

									end
									else
									if((r_sys_run_step==8'h6e)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1692[14:0] );

									end
									else
									if((r_sys_run_step==8'h2f)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1314[14:0] );

									end
									else
									if((r_sys_run_step==8'h29)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1278[14:0] );

									end
									else
									if((r_sys_run_step==8'h59)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp1566[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h23) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h86)) begin
										r_sub05_u_datain <= w_sys_tmp1046;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h23) || (r_sys_run_step==8'h26) || (r_sys_run_step==8'h29) || (r_sys_run_step==8'h2c) || (r_sys_run_step==8'h2f) || (r_sys_run_step==8'h32) || (r_sys_run_step==8'h35) || (r_sys_run_step==8'h38) || (r_sys_run_step==8'h3b) || (r_sys_run_step==8'h3e) || (r_sys_run_step==8'h41) || (r_sys_run_step==8'h44) || (r_sys_run_step==8'h47) || (r_sys_run_step==8'h4a) || (r_sys_run_step==8'h4d) || (r_sys_run_step==8'h50) || (r_sys_run_step==8'h53) || (r_sys_run_step==8'h56) || (r_sys_run_step==8'h59) || (r_sys_run_step==8'h5c) || (r_sys_run_step==8'h5f) || (r_sys_run_step==8'h62) || (r_sys_run_step==8'h65) || (r_sys_run_step==8'h68) || (r_sys_run_step==8'h6b) || (r_sys_run_step==8'h6e) || (r_sys_run_step==8'h71) || (r_sys_run_step==8'h74) || (r_sys_run_step==8'h77) || (r_sys_run_step==8'h7a) || (r_sys_run_step==8'h7d) || (r_sys_run_step==8'h80) || (r_sys_run_step==8'h83) || (r_sys_run_step==8'h86)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2778[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2958[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2988[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3153[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2838[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3183[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3003[14:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2718[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2943[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3108[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2868[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2823[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2898[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2853[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3063[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2913[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3123[14:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2733[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2763[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2808[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3168[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2883[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3033[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3138[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3078[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2748[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2973[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2793[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2928[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3048[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3093[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp3018[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1f)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1188[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1140[14:0] );

									end
									else
									if((r_sys_run_step==8'h2)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1044[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1056[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1050[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1176[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1086[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1134[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1110[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1122[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1068[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1164[14:0] );

									end
									else
									if((r_sys_run_step==8'h21)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1230[14:0] );

									end
									else
									if((r_sys_run_step==8'h1f)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1218[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1116[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1194[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1158[14:0] );

									end
									else
									if((r_sys_run_step==8'h22)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1236[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1200[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1146[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1182[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1206[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1152[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1098[14:0] );

									end
									else
									if((r_sys_run_step==8'h20)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1224[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1074[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1128[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1212[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1092[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1170[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1080[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1062[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp1104[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h22)) begin
										r_sub04_u_datain <= w_sys_tmp1046;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h2<=r_sys_run_step && r_sys_run_step<=8'h22)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2544[14:0] );

									end
									else
									if((r_sys_run_step==8'h16)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2664[14:0] );

									end
									else
									if((r_sys_run_step==8'h18)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2676[14:0] );

									end
									else
									if((r_sys_run_step==8'h9)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2586[14:0] );

									end
									else
									if((r_sys_run_step==8'hc)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2604[14:0] );

									end
									else
									if((r_sys_run_step==8'h4)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2556[14:0] );

									end
									else
									if((r_sys_run_step==8'h15)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2658[14:0] );

									end
									else
									if((r_sys_run_step==8'h1e)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2712[14:0] );

									end
									else
									if((r_sys_run_step==8'h19)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2682[14:0] );

									end
									else
									if((r_sys_run_step==8'h1c)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2700[14:0] );

									end
									else
									if((r_sys_run_step==8'h1a)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2688[14:0] );

									end
									else
									if((r_sys_run_step==8'hd)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2610[14:0] );

									end
									else
									if((r_sys_run_step==8'h7)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2574[14:0] );

									end
									else
									if((r_sys_run_step==8'h17)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2670[14:0] );

									end
									else
									if((r_sys_run_step==8'h13)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2646[14:0] );

									end
									else
									if((r_sys_run_step==8'hb)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2598[14:0] );

									end
									else
									if((r_sys_run_step==8'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2550[14:0] );

									end
									else
									if((r_sys_run_step==8'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2568[14:0] );

									end
									else
									if((r_sys_run_step==8'h1b)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2694[14:0] );

									end
									else
									if((r_sys_run_step==8'h10)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2628[14:0] );

									end
									else
									if((r_sys_run_step==8'h14)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2652[14:0] );

									end
									else
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2532[14:0] );

									end
									else
									if((r_sys_run_step==8'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2538[14:0] );

									end
									else
									if((r_sys_run_step==8'he)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2616[14:0] );

									end
									else
									if((r_sys_run_step==8'h12)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2640[14:0] );

									end
									else
									if((r_sys_run_step==8'h11)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2634[14:0] );

									end
									else
									if((r_sys_run_step==8'h8)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2580[14:0] );

									end
									else
									if((r_sys_run_step==8'hf)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2622[14:0] );

									end
									else
									if((r_sys_run_step==8'h1d)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2706[14:0] );

									end
									else
									if((r_sys_run_step==8'ha)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2592[14:0] );

									end
									else
									if((r_sys_run_step==8'h5)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2562[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h25: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==8'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((8'h0<=r_sys_run_step && r_sys_run_step<=8'h1e)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						6'h37: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h21)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h21)) begin
										r_sys_tmp0_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						6'h35: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp0_float <= w_sys_tmp3198;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h21)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h21)) begin
										r_sys_tmp1_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_tmp2_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_tmp2_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_tmp3_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_tmp3_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_tmp4_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h20)) begin
										r_sys_tmp4_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1f)) begin
										r_sys_tmp5_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1f)) begin
										r_sys_tmp5_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1f)) begin
										r_sys_tmp6_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1f)) begin
										r_sys_tmp6_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1f)) begin
										r_sys_tmp7_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1f)) begin
										r_sys_tmp7_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_tmp8_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_tmp8_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_tmp9_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_tmp9_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_tmp10_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1e)) begin
										r_sys_tmp10_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1d)) begin
										r_sys_tmp11_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1d)) begin
										r_sys_tmp11_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1d)) begin
										r_sys_tmp12_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1d)) begin
										r_sys_tmp12_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1d)) begin
										r_sys_tmp13_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1d)) begin
										r_sys_tmp13_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1c)) begin
										r_sys_tmp14_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1c)) begin
										r_sys_tmp14_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1c)) begin
										r_sys_tmp15_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1c)) begin
										r_sys_tmp15_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1c)) begin
										r_sys_tmp16_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sys_tmp16_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sys_tmp17_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1c)) begin
										r_sys_tmp17_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sys_tmp18_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sys_tmp18_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sys_tmp19_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1b)) begin
										r_sys_tmp19_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sys_tmp20_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sys_tmp20_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sys_tmp21_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sys_tmp21_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sys_tmp22_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_sys_tmp22_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_sys_tmp23_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h1a)) begin
										r_sys_tmp23_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_sys_tmp24_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_sys_tmp24_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_sys_tmp25_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h19)) begin
										r_sys_tmp25_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sys_tmp26_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sys_tmp26_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sys_tmp27_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sys_tmp27_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sys_tmp28_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h17)) begin
										r_sys_tmp28_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h17)) begin
										r_sys_tmp29_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h18)) begin
										r_sys_tmp29_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h17)) begin
										r_sys_tmp30_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h17)) begin
										r_sys_tmp30_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h17)) begin
										r_sys_tmp31_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h17)) begin
										r_sys_tmp31_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp32_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp32_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp33_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sys_tmp33_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp34_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp34_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sys_tmp35_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h16)) begin
										r_sys_tmp35_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sys_tmp36_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_tmp36_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sys_tmp37_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_tmp37_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_tmp38_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sys_tmp38_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_tmp39_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h15)) begin
										r_sys_tmp39_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_tmp40_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h13)) begin
										r_sys_tmp40_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h13)) begin
										r_sys_tmp41_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h13)) begin
										r_sys_tmp41_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h13)) begin
										r_sys_tmp42_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h14)) begin
										r_sys_tmp42_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h13)) begin
										r_sys_tmp43_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h13)) begin
										r_sys_tmp43_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_tmp44_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_tmp44_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_tmp45_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h11)) begin
										r_sys_tmp45_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_tmp46_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_tmp46_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h11)) begin
										r_sys_tmp47_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h12)) begin
										r_sys_tmp47_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h11)) begin
										r_sys_tmp48_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h10)) begin
										r_sys_tmp48_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h11)) begin
										r_sys_tmp49_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h10)) begin
										r_sys_tmp49_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h10)) begin
										r_sys_tmp50_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h11)) begin
										r_sys_tmp50_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h10)) begin
										r_sys_tmp51_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h11)) begin
										r_sys_tmp51_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h10)) begin
										r_sys_tmp52_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hf)) begin
										r_sys_tmp52_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hf)) begin
										r_sys_tmp53_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hf)) begin
										r_sys_tmp53_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hf)) begin
										r_sys_tmp54_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hf)) begin
										r_sys_tmp54_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hf)) begin
										r_sys_tmp55_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h10)) begin
										r_sys_tmp55_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'he)) begin
										r_sys_tmp56_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_tmp56_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'he)) begin
										r_sys_tmp57_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'he)) begin
										r_sys_tmp57_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'he)) begin
										r_sys_tmp58_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'he)) begin
										r_sys_tmp58_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_tmp59_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'he)) begin
										r_sys_tmp59_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_tmp60_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_sys_tmp60_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_tmp61_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_sys_tmp61_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_sys_tmp62_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_tmp62_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_sys_tmp63_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hd)) begin
										r_sys_tmp63_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_sys_tmp64_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sys_tmp64_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hb)) begin
										r_sys_tmp65_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sys_tmp65_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hb)) begin
										r_sys_tmp66_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sys_tmp66_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hb)) begin
										r_sys_tmp67_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h9)) begin
										r_sys_tmp67_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sys_tmp68_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hc)) begin
										r_sys_tmp68_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sys_tmp69_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hb)) begin
										r_sys_tmp69_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'ha)) begin
										r_sys_tmp70_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hb)) begin
										r_sys_tmp70_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h9)) begin
										r_sys_tmp71_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'hb)) begin
										r_sys_tmp71_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h9)) begin
										r_sys_tmp72_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp72_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h9)) begin
										r_sys_tmp73_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp73_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp74_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp74_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp75_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp75_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp76_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h9)) begin
										r_sys_tmp76_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp77_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h9)) begin
										r_sys_tmp77_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp78_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp78_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h7)) begin
										r_sys_tmp79_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h8)) begin
										r_sys_tmp79_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp80_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp80_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp81_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp81_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp82_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp82_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp83_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp83_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp84_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp84_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp85_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp85_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp86_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h5)) begin
										r_sys_tmp86_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp87_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h6)) begin
										r_sys_tmp87_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp88_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp88_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp89_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp89_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp90_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp90_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp91_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp91_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp92_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h3)) begin
										r_sys_tmp92_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2)) begin
										r_sys_tmp93_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h4)) begin
										r_sys_tmp93_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						6'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h21)) begin
										r_sys_tmp94_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						6'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==8'h2) || (r_sys_run_step==8'h21)) begin
										r_sys_tmp94_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
