/*
TimeStamp:	2016/10/20		16:0
*/


module sub07(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy,	
	input  signed  [14:0] i_fld_T_0_addr_0,	
	input          [31:0] i_fld_T_0_datain_0,	
	output         [31:0] o_fld_T_0_dataout_0,	
	input                 i_fld_T_0_r_w_0,	
	input  signed  [14:0] i_fld_V_1_addr_0,	
	input          [31:0] i_fld_V_1_datain_0,	
	output         [31:0] o_fld_V_1_dataout_0,	
	input                 i_fld_V_1_r_w_0,	
	input  signed  [14:0] i_fld_U_2_addr_0,	
	input          [31:0] i_fld_U_2_datain_0,	
	output         [31:0] o_fld_U_2_dataout_0,	
	input                 i_fld_U_2_r_w_0,	
	input  signed  [14:0] i_fld_result_3_addr_0,	
	input          [31:0] i_fld_result_3_datain_0,	
	output         [31:0] o_fld_result_3_dataout_0,	
	input                 i_fld_result_3_r_w_0	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 4:0] r_sys_run_phase;
	reg         [ 1:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 1:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [14:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [14:0] w_fld_V_1_addr_0;
	wire        [31:0] w_fld_V_1_datain_0;
	wire        [31:0] w_fld_V_1_dataout_0;
	wire               w_fld_V_1_r_w_0;
	wire               w_fld_V_1_ce_0;
	reg  signed [14:0] r_fld_V_1_addr_1;
	reg         [31:0] r_fld_V_1_datain_1;
	wire        [31:0] w_fld_V_1_dataout_1;
	reg                r_fld_V_1_r_w_1;
	wire               w_fld_V_1_ce_1;
	wire signed [14:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [14:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [14:0] w_fld_result_3_addr_0;
	wire        [31:0] w_fld_result_3_datain_0;
	wire        [31:0] w_fld_result_3_dataout_0;
	wire               w_fld_result_3_r_w_0;
	wire               w_fld_result_3_ce_0;
	reg  signed [14:0] r_fld_result_3_addr_1;
	reg         [31:0] r_fld_result_3_datain_1;
	wire        [31:0] w_fld_result_3_dataout_1;
	reg                r_fld_result_3_r_w_1;
	wire               w_fld_result_3_ce_1;
	reg  signed [31:0] r_run_k_4;
	reg  signed [31:0] r_run_j_5;
	reg  signed [31:0] r_run_kx_6;
	reg  signed [31:0] r_run_ky_7;
	reg  signed [31:0] r_run_mx_8;
	reg  signed [31:0] r_run_my_9;
	reg         [31:0] r_run_dt_10;
	reg         [31:0] r_run_dx_11;
	reg         [31:0] r_run_dy_12;
	reg         [31:0] r_run_r1_13;
	reg         [31:0] r_run_r2_14;
	reg         [31:0] r_run_r3_15;
	reg         [31:0] r_run_r4_16;
	reg         [31:0] r_run_YY_17;
	reg  signed [31:0] r_run_copy0_j_18;
	reg  signed [31:0] r_run_copy0_j_19;
	reg  signed [31:0] r_run_copy1_j_20;
	reg  signed [31:0] r_run_copy2_j_21;
	reg  signed [31:0] r_run_copy3_j_22;
	reg  signed [31:0] r_run_copy4_j_23;
	reg  signed [31:0] r_run_copy5_j_24;
	reg  signed [31:0] r_run_copy6_j_25;
	reg  signed [31:0] r_run_copy7_j_26;
	reg  signed [31:0] r_run_copy8_j_27;
	reg  signed [31:0] r_run_copy9_j_28;
	reg  signed [31:0] r_run_copy10_j_29;
	reg  signed [31:0] r_run_copy11_j_30;
	reg  signed [31:0] r_run_copy12_j_31;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire               w_sys_tmp12;
	wire               w_sys_tmp13;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp17;
	wire        [31:0] w_sys_tmp18;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire        [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire signed [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp26;
	wire signed [31:0] w_sys_tmp28;
	wire               w_sys_tmp29;
	wire               w_sys_tmp30;
	wire signed [31:0] w_sys_tmp31;
	wire signed [31:0] w_sys_tmp34;
	wire signed [31:0] w_sys_tmp35;
	wire signed [31:0] w_sys_tmp36;
	wire        [31:0] w_sys_tmp37;
	wire signed [31:0] w_sys_tmp39;
	wire signed [31:0] w_sys_tmp40;
	wire signed [31:0] w_sys_tmp43;
	wire signed [31:0] w_sys_tmp44;
	wire signed [31:0] w_sys_tmp93;
	wire               w_sys_tmp94;
	wire               w_sys_tmp95;
	wire signed [31:0] w_sys_tmp96;
	wire signed [31:0] w_sys_tmp97;
	wire signed [31:0] w_sys_tmp98;
	wire               w_sys_tmp99;
	wire               w_sys_tmp100;
	wire signed [31:0] w_sys_tmp101;
	wire signed [31:0] w_sys_tmp104;
	wire signed [31:0] w_sys_tmp105;
	wire signed [31:0] w_sys_tmp106;
	wire        [31:0] w_sys_tmp107;
	wire signed [31:0] w_sys_tmp108;
	wire signed [31:0] w_sys_tmp109;
	wire        [31:0] w_sys_tmp111;
	wire        [31:0] w_sys_tmp112;
	wire signed [31:0] w_sys_tmp113;
	wire signed [31:0] w_sys_tmp114;
	wire signed [31:0] w_sys_tmp117;
	wire signed [31:0] w_sys_tmp118;
	wire signed [31:0] w_sys_tmp119;
	wire        [31:0] w_sys_tmp121;
	wire signed [31:0] w_sys_tmp122;
	wire signed [31:0] w_sys_tmp123;
	wire signed [31:0] w_sys_tmp124;
	wire signed [31:0] w_sys_tmp127;
	wire signed [31:0] w_sys_tmp128;
	wire signed [31:0] w_sys_tmp130;
	wire signed [31:0] w_sys_tmp131;
	wire signed [31:0] w_sys_tmp132;
	wire signed [31:0] w_sys_tmp135;
	wire signed [31:0] w_sys_tmp136;
	wire signed [31:0] w_sys_tmp137;
	wire signed [31:0] w_sys_tmp140;
	wire signed [31:0] w_sys_tmp141;
	wire signed [31:0] w_sys_tmp142;
	wire        [31:0] w_sys_tmp145;
	wire signed [31:0] w_sys_tmp147;
	wire signed [31:0] w_sys_tmp148;
	wire signed [31:0] w_sys_tmp150;
	wire signed [31:0] w_sys_tmp151;
	wire signed [31:0] w_sys_tmp152;
	wire signed [31:0] w_sys_tmp156;
	wire signed [31:0] w_sys_tmp157;
	wire signed [31:0] w_sys_tmp158;
	wire signed [31:0] w_sys_tmp163;
	wire signed [31:0] w_sys_tmp164;
	wire signed [31:0] w_sys_tmp166;
	wire signed [31:0] w_sys_tmp167;
	wire signed [31:0] w_sys_tmp168;
	wire signed [31:0] w_sys_tmp170;
	wire signed [31:0] w_sys_tmp171;
	wire signed [31:0] w_sys_tmp172;
	wire signed [31:0] w_sys_tmp173;
	wire signed [31:0] w_sys_tmp174;
	wire signed [31:0] w_sys_tmp176;
	wire signed [31:0] w_sys_tmp177;
	wire signed [31:0] w_sys_tmp178;
	wire signed [31:0] w_sys_tmp179;
	wire signed [31:0] w_sys_tmp181;
	wire signed [31:0] w_sys_tmp182;
	wire signed [31:0] w_sys_tmp183;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 2'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign o_fld_T_0_dataout_0 = w_fld_T_0_dataout_0;
	assign w_fld_T_0_addr_0 = i_fld_T_0_addr_0;
	assign w_fld_T_0_datain_0 = i_fld_T_0_datain_0;
	assign w_fld_T_0_r_w_0 = i_fld_T_0_r_w_0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign o_fld_V_1_dataout_0 = w_fld_V_1_dataout_0;
	assign w_fld_V_1_addr_0 = i_fld_V_1_addr_0;
	assign w_fld_V_1_datain_0 = i_fld_V_1_datain_0;
	assign w_fld_V_1_r_w_0 = i_fld_V_1_r_w_0;
	assign w_fld_V_1_ce_0 = w_sys_ce;
	assign w_fld_V_1_ce_1 = w_sys_ce;
	assign o_fld_U_2_dataout_0 = w_fld_U_2_dataout_0;
	assign w_fld_U_2_addr_0 = i_fld_U_2_addr_0;
	assign w_fld_U_2_datain_0 = i_fld_U_2_datain_0;
	assign w_fld_U_2_r_w_0 = i_fld_U_2_r_w_0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign o_fld_result_3_dataout_0 = w_fld_result_3_dataout_0;
	assign w_fld_result_3_addr_0 = i_fld_result_3_addr_0;
	assign w_fld_result_3_datain_0 = i_fld_result_3_datain_0;
	assign w_fld_result_3_r_w_0 = i_fld_result_3_r_w_0;
	assign w_fld_result_3_ce_0 = w_sys_ce;
	assign w_fld_result_3_ce_1 = w_sys_ce;
	assign w_sys_tmp1 = 32'sh00000080;
	assign w_sys_tmp3 = 32'sh00000081;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'h3d000000;
	assign w_sys_tmp7 = 32'h3c000000;
	assign w_sys_tmp8 = 32'h3c03126f;
	assign w_sys_tmp9 = 32'h3d03126f;
	assign w_sys_tmp10 = 32'h3f03126f;
	assign w_sys_tmp11 = 32'h4103126f;
	assign w_sys_tmp12 = ( !w_sys_tmp13 );
	assign w_sys_tmp13 = (r_run_my_9 < r_run_k_4);
	assign w_sys_tmp16 = (w_sys_tmp17 + r_run_k_4);
	assign w_sys_tmp17 = 32'sh00000081;
	assign w_sys_tmp18 = 32'h0;
	assign w_sys_tmp20 = (w_sys_tmp21 + r_run_k_4);
	assign w_sys_tmp21 = (r_run_mx_8 * w_sys_tmp17);
	assign w_sys_tmp23 = w_fld_T_0_dataout_1;
	assign w_sys_tmp24 = (w_sys_tmp25 + r_run_k_4);
	assign w_sys_tmp25 = (w_sys_tmp26 * w_sys_tmp17);
	assign w_sys_tmp26 = (r_run_mx_8 - w_sys_intOne);
	assign w_sys_tmp28 = (r_run_k_4 + w_sys_intOne);
	assign w_sys_tmp29 = ( !w_sys_tmp30 );
	assign w_sys_tmp30 = (w_sys_tmp31 < r_run_j_5);
	assign w_sys_tmp31 = 32'sh00000022;
	assign w_sys_tmp34 = (w_sys_tmp35 + w_sys_intOne);
	assign w_sys_tmp35 = (r_run_j_5 * w_sys_tmp36);
	assign w_sys_tmp36 = 32'sh00000081;
	assign w_sys_tmp37 = 32'h0;
	assign w_sys_tmp39 = (w_sys_tmp40 + r_run_my_9);
	assign w_sys_tmp40 = (r_run_copy0_j_18 * w_sys_tmp36);
	assign w_sys_tmp43 = (r_run_copy0_j_18 + w_sys_intOne);
	assign w_sys_tmp44 = (r_run_j_5 + w_sys_intOne);
	assign w_sys_tmp93 = 32'sh00000021;
	assign w_sys_tmp94 = ( !w_sys_tmp95 );
	assign w_sys_tmp95 = (w_sys_tmp96 < r_run_k_4);
	assign w_sys_tmp96 = 32'sh00000040;
	assign w_sys_tmp97 = (r_run_k_4 + w_sys_intOne);
	assign w_sys_tmp98 = 32'sh00000002;
	assign w_sys_tmp99 = ( !w_sys_tmp100 );
	assign w_sys_tmp100 = (w_sys_tmp101 < r_run_j_5);
	assign w_sys_tmp101 = 32'sh00000021;
	assign w_sys_tmp104 = (w_sys_tmp105 + r_run_k_4);
	assign w_sys_tmp105 = (r_run_j_5 * w_sys_tmp106);
	assign w_sys_tmp106 = 32'sh00000081;
	assign w_sys_tmp107 = w_ip_AddFloat_result_0;
	assign w_sys_tmp108 = (w_sys_tmp109 + r_run_k_4);
	assign w_sys_tmp109 = (r_run_copy12_j_31 * w_sys_tmp106);
	assign w_sys_tmp111 = w_ip_MultFloat_product_0;
	assign w_sys_tmp112 = w_fld_U_2_dataout_1;
	assign w_sys_tmp113 = (w_sys_tmp114 + r_run_k_4);
	assign w_sys_tmp114 = (r_run_copy11_j_30 * w_sys_tmp106);
	assign w_sys_tmp117 = (w_sys_tmp118 + r_run_k_4);
	assign w_sys_tmp118 = (w_sys_tmp119 * w_sys_tmp106);
	assign w_sys_tmp119 = (r_run_copy10_j_29 + w_sys_intOne);
	assign w_sys_tmp121 = w_fld_T_0_dataout_1;
	assign w_sys_tmp122 = (w_sys_tmp123 + r_run_k_4);
	assign w_sys_tmp123 = (w_sys_tmp124 * w_sys_tmp106);
	assign w_sys_tmp124 = (r_run_copy9_j_28 - w_sys_intOne);
	assign w_sys_tmp127 = (w_sys_tmp128 + r_run_k_4);
	assign w_sys_tmp128 = (r_run_copy8_j_27 * w_sys_tmp106);
	assign w_sys_tmp130 = (w_sys_tmp131 + w_sys_intOne);
	assign w_sys_tmp131 = (w_sys_tmp132 + r_run_k_4);
	assign w_sys_tmp132 = (r_run_copy7_j_26 * w_sys_tmp106);
	assign w_sys_tmp135 = (w_sys_tmp136 - w_sys_intOne);
	assign w_sys_tmp136 = (w_sys_tmp137 + r_run_k_4);
	assign w_sys_tmp137 = (r_run_copy6_j_25 * w_sys_tmp106);
	assign w_sys_tmp140 = (w_sys_tmp141 + r_run_k_4);
	assign w_sys_tmp141 = (w_sys_tmp142 * w_sys_tmp106);
	assign w_sys_tmp142 = (r_run_copy5_j_24 + w_sys_intOne);
	assign w_sys_tmp145 = 32'h40000000;
	assign w_sys_tmp147 = (w_sys_tmp148 + r_run_k_4);
	assign w_sys_tmp148 = (r_run_copy4_j_23 * w_sys_tmp106);
	assign w_sys_tmp150 = (w_sys_tmp151 + r_run_k_4);
	assign w_sys_tmp151 = (w_sys_tmp152 * w_sys_tmp106);
	assign w_sys_tmp152 = (r_run_copy3_j_22 - w_sys_intOne);
	assign w_sys_tmp156 = (w_sys_tmp157 + w_sys_intOne);
	assign w_sys_tmp157 = (w_sys_tmp158 + r_run_k_4);
	assign w_sys_tmp158 = (r_run_copy2_j_21 * w_sys_tmp106);
	assign w_sys_tmp163 = (w_sys_tmp164 + r_run_k_4);
	assign w_sys_tmp164 = (r_run_copy1_j_20 * w_sys_tmp106);
	assign w_sys_tmp166 = (w_sys_tmp167 - w_sys_intOne);
	assign w_sys_tmp167 = (w_sys_tmp168 + r_run_k_4);
	assign w_sys_tmp168 = (r_run_copy0_j_19 * w_sys_tmp106);
	assign w_sys_tmp170 = (r_run_copy0_j_19 + w_sys_intOne);
	assign w_sys_tmp171 = (r_run_copy1_j_20 + w_sys_intOne);
	assign w_sys_tmp172 = (r_run_copy2_j_21 + w_sys_intOne);
	assign w_sys_tmp173 = (r_run_copy3_j_22 + w_sys_intOne);
	assign w_sys_tmp174 = (r_run_copy4_j_23 + w_sys_intOne);
	assign w_sys_tmp176 = (r_run_copy6_j_25 + w_sys_intOne);
	assign w_sys_tmp177 = (r_run_copy7_j_26 + w_sys_intOne);
	assign w_sys_tmp178 = (r_run_copy8_j_27 + w_sys_intOne);
	assign w_sys_tmp179 = (r_run_copy9_j_28 + w_sys_intOne);
	assign w_sys_tmp181 = (r_run_copy11_j_30 + w_sys_intOne);
	assign w_sys_tmp182 = (r_run_copy12_j_31 + w_sys_intOne);
	assign w_sys_tmp183 = (r_run_j_5 + w_sys_intOne);


	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_V_1(
			.clk (clock),
			.ce_0 (w_fld_V_1_ce_0),
			.addr_0 (w_fld_V_1_addr_0),
			.datain_0 (w_fld_V_1_datain_0),
			.dataout_0 (w_fld_V_1_dataout_0),
			.r_w_0 (w_fld_V_1_r_w_0),
			.ce_1 (w_fld_V_1_ce_1),
			.addr_1 (r_fld_V_1_addr_1),
			.datain_1 (r_fld_V_1_datain_1),
			.dataout_1 (w_fld_V_1_dataout_1),
			.r_w_1 (r_fld_V_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_result_3(
			.clk (clock),
			.ce_0 (w_fld_result_3_ce_0),
			.addr_0 (w_fld_result_3_addr_0),
			.datain_0 (w_fld_result_3_datain_0),
			.dataout_0 (w_fld_result_3_dataout_0),
			.r_w_0 (w_fld_result_3_r_w_0),
			.ce_1 (w_fld_result_3_ce_1),
			.addr_1 (r_fld_result_3_addr_1),
			.datain_1 (r_fld_result_3_datain_1),
			.dataout_1 (w_fld_result_3_dataout_1),
			.r_w_1 (r_fld_result_3_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h2c) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h3b)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h3c)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h3a)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'h12) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h3e) || (r_sys_run_step==7'h3f) || (r_sys_run_step==7'h41) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h4d)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp107;

									end
									else
									if((r_sys_run_step==7'h14) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h48)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h39)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp12_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp121[31], w_sys_tmp121[30:0] };

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp121[31], w_sys_tmp121[30:0] };

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp121[31], w_sys_tmp121[30:0] };

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp7_float[31], r_sys_tmp7_float[30:0] };

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp121[31], w_sys_tmp121[30:0] };

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h15) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h36) || (r_sys_run_step==7'h41)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp121[31], w_sys_tmp121[30:0] };

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp121[31], w_sys_tmp121[30:0] };

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp121[31], w_sys_tmp121[30:0] };

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp11_float[31], r_sys_tmp11_float[30:0] };

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp121[31], w_sys_tmp121[30:0] };

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp7_float[31], r_sys_tmp7_float[30:0] };

									end
									else
									if((r_sys_run_step==7'h37) || (r_sys_run_step==7'h40)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp121[31], w_sys_tmp121[30:0] };

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp121[31], w_sys_tmp121[30:0] };

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_ip_AddFloat_portB_0 <= { ~r_sys_tmp11_float[31], r_sys_tmp11_float[30:0] };

									end
									else
									if((r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2a)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h12) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h33) || (r_sys_run_step==7'h3e)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h48)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp111;

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp111[31], w_sys_tmp111[30:0] };

									end
									else
									if((r_sys_run_step==7'h2c) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h45) || (r_sys_run_step==7'h4d)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp11_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h2a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'hf) || (r_sys_run_step==7'h17)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h8) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h37)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp145;

									end
									else
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'he)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r2_14;

									end
									else
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h43)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r3_15;

									end
									else
									if((r_sys_run_step==7'h1a) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h46)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r4_16;

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp7_float;

									end
									else
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_r1_13;

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h1f)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp11_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hc)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp9_float;

									end
									else
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp112;

									end
									else
									if((r_sys_run_step==7'h8) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h34) || (r_sys_run_step==7'h37)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp121;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h30) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h3b) || (r_sys_run_step==7'h43) || (r_sys_run_step==7'h46)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp107;

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h39)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp11_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						5'h1b: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h0: begin
							r_sys_run_phase <= 5'h2;
						end

						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 5'h4;

									end
								end

							endcase
						end

						5'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 5'h5;

									end
								end

							endcase
						end

						5'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12) ? 5'h8 : 5'ha);

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_run_phase <= 5'h5;

									end
								end

							endcase
						end

						5'ha: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 5'hb;

									end
								end

							endcase
						end

						5'hb: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp29) ? 5'he : 5'h10);

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_run_phase <= 5'hb;

									end
								end

							endcase
						end

						5'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 5'h11;

									end
								end

							endcase
						end

						5'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp94) ? 5'h15 : 5'h1b);

									end
								end

							endcase
						end

						5'h12: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 5'h11;

									end
								end

							endcase
						end

						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 5'h16;

									end
								end

							endcase
						end

						5'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp99) ? 5'h19 : 5'h12);

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h52)) begin
										r_sys_run_phase <= 5'h16;

									end
								end

							endcase
						end

						5'h1b: begin
							r_sys_run_phase <= 5'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'hb: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h12: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h52)) begin
										r_sys_run_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'h5: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'hb: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'h11: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'h12: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'h16: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h51)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h52)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						5'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						5'h1b: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp24[14:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp20[14:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp16[14:0] );

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp39[14:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h2) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp34[14:0] );

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h35)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp163[14:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h36)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp166[14:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp108[14:0] );

									end
									else
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp135[14:0] );

									end
									else
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp130[14:0] );

									end
									else
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp122[14:0] );

									end
									else
									if((r_sys_run_step==7'h8) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp156[14:0] );

									end
									else
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp140[14:0] );

									end
									else
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp150[14:0] );

									end
									else
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp117[14:0] );

									end
									else
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp147[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp23;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp37;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h3)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h36)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						5'h1b: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_1_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4)) begin
										r_fld_V_1_addr_1 <= $signed( w_sys_tmp127[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4)) begin
										r_fld_V_1_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						5'h1b: begin
							r_fld_V_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp113[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						5'h1b: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_result_3_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h31) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h52)) begin
										r_fld_result_3_addr_1 <= $signed( w_sys_tmp104[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h31) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h52)) begin
										r_fld_result_3_datain_1 <= w_sys_tmp107;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_result_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h31) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h52)) begin
										r_fld_result_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						5'h1b: begin
							r_fld_result_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h4: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_4 <= w_sys_intOne;

									end
								end

							endcase
						end

						5'h8: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_run_k_4 <= w_sys_tmp28;

									end
								end

							endcase
						end

						5'h10: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_4 <= w_sys_tmp93;

									end
								end

							endcase
						end

						5'h12: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_4 <= w_sys_tmp97;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'ha: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_5 <= w_sys_intOne;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h2) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h8)) begin
										r_run_j_5 <= w_sys_tmp44;

									end
								end

							endcase
						end

						5'h15: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_5 <= w_sys_tmp98;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h31) || (r_sys_run_step==7'h3c) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h4a) || (r_sys_run_step==7'h52)) begin
										r_run_j_5 <= w_sys_tmp183;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_kx_6 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_ky_7 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_mx_8 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_my_9 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dt_10 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dx_11 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dy_12 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r1_13 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r2_14 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r3_15 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h2: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r4_16 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'ha: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_18 <= r_run_j_5;

									end
								end

							endcase
						end

						5'he: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9)) begin
										r_run_copy0_j_18 <= w_sys_tmp43;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_19 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h36)) begin
										r_run_copy0_j_19 <= w_sys_tmp170;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_20 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h35)) begin
										r_run_copy1_j_20 <= w_sys_tmp171;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_21 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h8) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h1e) || (r_sys_run_step==7'h29) || (r_sys_run_step==7'h34)) begin
										r_run_copy2_j_21 <= w_sys_tmp172;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy3_j_22 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h33)) begin
										r_run_copy3_j_22 <= w_sys_tmp173;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy4_j_23 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h6) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h32)) begin
										r_run_copy4_j_23 <= w_sys_tmp174;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy5_j_24 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h5) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h31)) begin
										r_run_copy5_j_24 <= w_sys_tmp142;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy6_j_25 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h4) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1a) || (r_sys_run_step==7'h25) || (r_sys_run_step==7'h30)) begin
										r_run_copy6_j_25 <= w_sys_tmp176;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy7_j_26 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h2f)) begin
										r_run_copy7_j_26 <= w_sys_tmp177;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy8_j_27 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4)) begin
										r_run_copy8_j_27 <= w_sys_tmp178;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy9_j_28 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2e)) begin
										r_run_copy9_j_28 <= w_sys_tmp179;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy10_j_29 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'hc) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2d)) begin
										r_run_copy10_j_29 <= w_sys_tmp119;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy11_j_30 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h4)) begin
										r_run_copy11_j_30 <= w_sys_tmp181;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h15: begin

							case(r_sys_run_stage) 
								2'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy12_j_31 <= r_run_j_5;

									end
								end

							endcase
						end

						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h2c)) begin
										r_run_copy12_j_31 <= w_sys_tmp182;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h12)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp1_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h33)) begin
										r_sys_tmp2_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h13)) begin
										r_sys_tmp3_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp3_float <= w_fld_V_1_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'hf) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h28)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h20) || (r_sys_run_step==7'h2b) || (r_sys_run_step==7'h36)) begin
										r_sys_tmp5_float <= w_fld_T_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h9) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h35)) begin
										r_sys_tmp6_float <= w_fld_T_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h8) || (r_sys_run_step==7'h1c) || (r_sys_run_step==7'h27) || (r_sys_run_step==7'h2a) || (r_sys_run_step==7'h3e)) begin
										r_sys_tmp7_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h11)) begin
										r_sys_tmp8_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp8_float <= w_fld_V_1_dataout_1;

									end
									else
									if((r_sys_run_step==7'h24) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h3a)) begin
										r_sys_tmp8_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h38)) begin
										r_sys_tmp9_float <= w_fld_T_0_dataout_1;

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp9_float <= w_fld_V_1_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h2) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h24) || (r_sys_run_step==7'h26) || (r_sys_run_step==7'h28) || (r_sys_run_step==7'h2e)) begin
										r_sys_tmp10_float <= w_fld_T_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'h1f) || (r_sys_run_step==7'h32) || (r_sys_run_step==7'h35) || (r_sys_run_step==7'h3d) || (r_sys_run_step==7'h40) || (r_sys_run_step==7'h4b)) begin
										r_sys_tmp11_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp11_float <= w_fld_V_1_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1b) || (r_sys_run_step==7'h1d) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2f) || (r_sys_run_step==7'h31) || (r_sys_run_step==7'h33)) begin
										r_sys_tmp12_float <= w_fld_T_0_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						5'h19: begin

							case(r_sys_run_stage) 
								2'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp13_float <= w_fld_V_1_dataout_1;

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h16) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h21) || (r_sys_run_step==7'h22) || (r_sys_run_step==7'h23) || (r_sys_run_step==7'h2c) || (r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2e) || (r_sys_run_step==7'h37) || (r_sys_run_step==7'h38) || (r_sys_run_step==7'h39) || (r_sys_run_step==7'h44)) begin
										r_sys_tmp13_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
