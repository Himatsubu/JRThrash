/*
TimeStamp:	2016/10/27		16:53
*/


module P3_2dim(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 9:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 5:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 5:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [14:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [14:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [14:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [14:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [14:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [14:0] w_fld_V_3_addr_0;
	wire        [31:0] w_fld_V_3_datain_0;
	wire        [31:0] w_fld_V_3_dataout_0;
	wire               w_fld_V_3_r_w_0;
	wire               w_fld_V_3_ce_0;
	reg  signed [14:0] r_fld_V_3_addr_1;
	reg         [31:0] r_fld_V_3_datain_1;
	wire        [31:0] w_fld_V_3_dataout_1;
	reg                r_fld_V_3_r_w_1;
	wire               w_fld_V_3_ce_1;
	reg  signed [31:0] r_run_k_36;
	reg  signed [31:0] r_run_j_37;
	reg  signed [31:0] r_run_n_38;
	reg  signed [31:0] r_run_mx_39;
	reg  signed [31:0] r_run_my_40;
	reg         [31:0] r_run_dt_41;
	reg         [31:0] r_run_dx_42;
	reg         [31:0] r_run_dy_43;
	reg         [31:0] r_run_r1_44;
	reg         [31:0] r_run_r2_45;
	reg         [31:0] r_run_r3_46;
	reg         [31:0] r_run_r4_47;
	reg         [31:0] r_run_YY_48;
	reg  signed [31:0] r_run_kx_49;
	reg  signed [31:0] r_run_ky_50;
	reg  signed [31:0] r_run_nlast_51;
	reg  signed [31:0] r_run_tmpj_52;
	reg  signed [31:0] r_run_copy0_j_53;
	reg  signed [31:0] r_run_copy1_j_54;
	reg  signed [31:0] r_run_copy2_j_55;
	reg  signed [31:0] r_run_copy0_j_56;
	reg  signed [31:0] r_run_copy1_j_57;
	reg  signed [31:0] r_run_copy2_j_58;
	reg  signed [31:0] r_run_copy3_j_59;
	reg  signed [31:0] r_run_copy4_j_60;
	reg  signed [31:0] r_run_copy0_j_61;
	reg  signed [31:0] r_run_copy1_j_62;
	reg  signed [31:0] r_run_copy2_j_63;
	reg  signed [31:0] r_run_copy3_j_64;
	reg  signed [31:0] r_run_copy4_j_65;
	reg  signed [31:0] r_run_copy0_j_66;
	reg  signed [31:0] r_run_copy1_j_67;
	reg  signed [31:0] r_run_copy2_j_68;
	reg  signed [31:0] r_run_copy3_j_69;
	reg  signed [31:0] r_run_copy4_j_70;
	reg  signed [31:0] r_run_copy0_j_71;
	reg  signed [31:0] r_run_copy1_j_72;
	reg  signed [31:0] r_run_copy2_j_73;
	reg  signed [31:0] r_run_copy3_j_74;
	reg  signed [31:0] r_run_copy4_j_75;
	reg  signed [31:0] r_run_copy0_j_76;
	reg  signed [31:0] r_run_copy1_j_77;
	reg  signed [31:0] r_run_copy2_j_78;
	reg  signed [31:0] r_run_copy3_j_79;
	reg  signed [31:0] r_run_copy4_j_80;
	reg  signed [31:0] r_run_copy0_j_81;
	reg  signed [31:0] r_run_copy1_j_82;
	reg  signed [31:0] r_run_copy2_j_83;
	reg  signed [31:0] r_run_copy3_j_84;
	reg  signed [31:0] r_run_copy4_j_85;
	reg  signed [31:0] r_run_copy0_j_86;
	reg  signed [31:0] r_run_copy1_j_87;
	reg  signed [31:0] r_run_copy2_j_88;
	reg  signed [31:0] r_run_copy3_j_89;
	reg  signed [31:0] r_run_copy4_j_90;
	reg  signed [31:0] r_run_copy0_j_91;
	reg  signed [31:0] r_run_copy1_j_92;
	reg  signed [31:0] r_run_copy2_j_93;
	reg  signed [31:0] r_run_copy3_j_94;
	reg  signed [31:0] r_run_copy4_j_95;
	reg  signed [31:0] r_run_copy0_j_96;
	reg  signed [31:0] r_run_copy1_j_97;
	reg  signed [31:0] r_run_copy2_j_98;
	reg  signed [31:0] r_run_copy3_j_99;
	reg  signed [31:0] r_run_copy4_j_100;
	reg  signed [31:0] r_run_copy0_j_101;
	reg  signed [31:0] r_run_copy1_j_102;
	reg  signed [31:0] r_run_copy2_j_103;
	reg  signed [31:0] r_run_copy3_j_104;
	reg  signed [31:0] r_run_copy4_j_105;
	reg  signed [31:0] r_run_copy0_j_106;
	reg  signed [31:0] r_run_copy1_j_107;
	reg  signed [31:0] r_run_copy2_j_108;
	reg  signed [31:0] r_run_copy3_j_109;
	reg  signed [31:0] r_run_copy4_j_110;
	reg  signed [31:0] r_run_copy0_j_111;
	reg  signed [31:0] r_run_copy1_j_112;
	reg  signed [31:0] r_run_copy2_j_113;
	reg  signed [31:0] r_run_copy3_j_114;
	reg  signed [31:0] r_run_copy4_j_115;
	reg  signed [31:0] r_run_copy0_j_116;
	reg  signed [31:0] r_run_copy1_j_117;
	reg  signed [31:0] r_run_copy2_j_118;
	reg  signed [31:0] r_run_copy3_j_119;
	reg  signed [31:0] r_run_copy4_j_120;
	reg  signed [31:0] r_run_copy0_j_121;
	reg  signed [31:0] r_run_copy1_j_122;
	reg  signed [31:0] r_run_copy2_j_123;
	reg  signed [31:0] r_run_copy3_j_124;
	reg  signed [31:0] r_run_copy4_j_125;
	reg  signed [31:0] r_run_copy0_j_126;
	reg  signed [31:0] r_run_copy1_j_127;
	reg  signed [31:0] r_run_copy2_j_128;
	reg  signed [31:0] r_run_copy3_j_129;
	reg  signed [31:0] r_run_copy4_j_130;
	reg  signed [31:0] r_run_copy0_j_131;
	reg  signed [31:0] r_run_copy1_j_132;
	reg  signed [31:0] r_run_copy2_j_133;
	reg  signed [31:0] r_run_copy3_j_134;
	reg  signed [31:0] r_run_copy4_j_135;
	reg  signed [31:0] r_run_copy0_j_136;
	reg  signed [31:0] r_run_copy1_j_137;
	reg  signed [31:0] r_run_copy2_j_138;
	reg  signed [31:0] r_run_copy3_j_139;
	reg  signed [31:0] r_run_copy4_j_140;
	reg  signed [31:0] r_run_copy0_j_141;
	reg  signed [31:0] r_run_copy1_j_142;
	reg  signed [31:0] r_run_copy2_j_143;
	reg  signed [31:0] r_run_copy3_j_144;
	reg  signed [31:0] r_run_copy4_j_145;
	reg  signed [31:0] r_run_copy0_j_146;
	reg  signed [31:0] r_run_copy1_j_147;
	reg  signed [31:0] r_run_copy2_j_148;
	reg  signed [31:0] r_run_copy3_j_149;
	reg  signed [31:0] r_run_copy4_j_150;
	reg  signed [31:0] r_run_copy0_j_151;
	reg  signed [31:0] r_run_copy1_j_152;
	reg  signed [31:0] r_run_copy2_j_153;
	reg  signed [31:0] r_run_copy3_j_154;
	reg  signed [31:0] r_run_copy4_j_155;
	reg  signed [31:0] r_run_copy0_j_156;
	reg  signed [31:0] r_run_copy1_j_157;
	reg  signed [31:0] r_run_copy2_j_158;
	reg  signed [31:0] r_run_copy3_j_159;
	reg  signed [31:0] r_run_copy4_j_160;
	reg  signed [31:0] r_run_copy0_j_161;
	reg  signed [31:0] r_run_copy1_j_162;
	reg  signed [31:0] r_run_copy2_j_163;
	reg  signed [31:0] r_run_copy3_j_164;
	reg  signed [31:0] r_run_copy4_j_165;
	reg  signed [31:0] r_run_copy0_j_166;
	reg  signed [31:0] r_run_copy1_j_167;
	reg  signed [31:0] r_run_copy2_j_168;
	reg  signed [31:0] r_run_copy3_j_169;
	reg  signed [31:0] r_run_copy4_j_170;
	reg  signed [31:0] r_run_copy0_j_171;
	reg  signed [31:0] r_run_copy1_j_172;
	reg  signed [31:0] r_run_copy2_j_173;
	reg  signed [31:0] r_run_copy3_j_174;
	reg  signed [31:0] r_run_copy4_j_175;
	reg  signed [31:0] r_run_copy0_j_176;
	reg  signed [31:0] r_run_copy1_j_177;
	reg  signed [31:0] r_run_copy2_j_178;
	reg  signed [31:0] r_run_copy3_j_179;
	reg  signed [31:0] r_run_copy4_j_180;
	reg  signed [31:0] r_run_copy0_j_181;
	reg  signed [31:0] r_run_copy1_j_182;
	reg  signed [31:0] r_run_copy2_j_183;
	reg  signed [31:0] r_run_copy3_j_184;
	reg  signed [31:0] r_run_copy4_j_185;
	reg  signed [31:0] r_run_copy0_j_186;
	reg  signed [31:0] r_run_copy1_j_187;
	reg  signed [31:0] r_run_copy2_j_188;
	reg  signed [31:0] r_run_copy3_j_189;
	reg  signed [31:0] r_run_copy4_j_190;
	reg  signed [31:0] r_run_copy0_j_191;
	reg  signed [31:0] r_run_copy1_j_192;
	reg  signed [31:0] r_run_copy2_j_193;
	reg  signed [31:0] r_run_copy3_j_194;
	reg  signed [31:0] r_run_copy4_j_195;
	reg  signed [31:0] r_run_copy0_j_196;
	reg  signed [31:0] r_run_copy1_j_197;
	reg  signed [31:0] r_run_copy2_j_198;
	reg  signed [31:0] r_run_copy3_j_199;
	reg  signed [31:0] r_run_copy4_j_200;
	reg  signed [31:0] r_run_copy0_j_201;
	reg  signed [31:0] r_run_copy1_j_202;
	reg  signed [31:0] r_run_copy2_j_203;
	reg  signed [31:0] r_run_copy3_j_204;
	reg  signed [31:0] r_run_copy4_j_205;
	reg  signed [31:0] r_run_copy0_j_206;
	reg  signed [31:0] r_run_copy1_j_207;
	reg  signed [31:0] r_run_copy2_j_208;
	reg  signed [31:0] r_run_copy3_j_209;
	reg  signed [31:0] r_run_copy4_j_210;
	reg  signed [31:0] r_run_copy0_j_211;
	reg  signed [31:0] r_run_copy1_j_212;
	reg  signed [31:0] r_run_copy2_j_213;
	reg  signed [31:0] r_run_copy3_j_214;
	reg  signed [31:0] r_run_copy4_j_215;
	reg  signed [31:0] r_run_copy0_j_216;
	reg  signed [31:0] r_run_copy1_j_217;
	reg  signed [31:0] r_run_copy2_j_218;
	reg  signed [31:0] r_run_copy3_j_219;
	reg  signed [31:0] r_run_copy4_j_220;
	reg  signed [31:0] r_run_copy5_j_221;
	reg  signed [31:0] r_run_copy6_j_222;
	reg  signed [31:0] r_run_copy7_j_223;
	reg  signed [31:0] r_run_copy8_j_224;
	reg  signed [31:0] r_run_copy9_j_225;
	reg  signed [31:0] r_run_copy10_j_226;
	reg  signed [31:0] r_run_copy0_j_227;
	reg  signed [31:0] r_run_copy1_j_228;
	reg  signed [31:0] r_run_copy2_j_229;
	reg  signed [31:0] r_run_copy3_j_230;
	reg  signed [31:0] r_run_copy4_j_231;
	reg  signed [31:0] r_run_copy5_j_232;
	reg  signed [31:0] r_run_copy6_j_233;
	reg  signed [31:0] r_run_copy7_j_234;
	reg  signed [31:0] r_run_copy8_j_235;
	reg  signed [31:0] r_run_copy9_j_236;
	reg  signed [31:0] r_run_copy10_j_237;
	reg  signed [31:0] r_run_copy0_j_238;
	reg  signed [31:0] r_run_copy1_j_239;
	reg  signed [31:0] r_run_copy2_j_240;
	reg  signed [31:0] r_run_copy3_j_241;
	reg  signed [31:0] r_run_copy4_j_242;
	reg  signed [31:0] r_run_copy5_j_243;
	reg  signed [31:0] r_run_copy6_j_244;
	reg  signed [31:0] r_run_copy7_j_245;
	reg  signed [31:0] r_run_copy8_j_246;
	reg  signed [31:0] r_run_copy9_j_247;
	reg  signed [31:0] r_run_copy10_j_248;
	reg  signed [31:0] r_run_copy0_j_249;
	reg  signed [31:0] r_run_copy1_j_250;
	reg  signed [31:0] r_run_copy2_j_251;
	reg  signed [31:0] r_run_copy3_j_252;
	reg  signed [31:0] r_run_copy4_j_253;
	reg  signed [31:0] r_run_copy5_j_254;
	reg  signed [31:0] r_run_copy6_j_255;
	reg  signed [31:0] r_run_copy7_j_256;
	reg  signed [31:0] r_run_copy8_j_257;
	reg  signed [31:0] r_run_copy9_j_258;
	reg  signed [31:0] r_run_copy10_j_259;
	reg  signed [31:0] r_run_copy0_j_260;
	reg  signed [31:0] r_run_copy1_j_261;
	reg  signed [31:0] r_run_copy2_j_262;
	reg  signed [31:0] r_run_copy3_j_263;
	reg  signed [31:0] r_run_copy4_j_264;
	reg  signed [31:0] r_run_copy5_j_265;
	reg  signed [31:0] r_run_copy6_j_266;
	reg  signed [31:0] r_run_copy7_j_267;
	reg  signed [31:0] r_run_copy8_j_268;
	reg  signed [31:0] r_run_copy9_j_269;
	reg  signed [31:0] r_run_copy10_j_270;
	reg  signed [31:0] r_run_copy0_j_271;
	reg  signed [31:0] r_run_copy1_j_272;
	reg  signed [31:0] r_run_copy2_j_273;
	reg  signed [31:0] r_run_copy3_j_274;
	reg  signed [31:0] r_run_copy4_j_275;
	reg  signed [31:0] r_run_copy5_j_276;
	reg  signed [31:0] r_run_copy6_j_277;
	reg  signed [31:0] r_run_copy7_j_278;
	reg  signed [31:0] r_run_copy8_j_279;
	reg  signed [31:0] r_run_copy9_j_280;
	reg  signed [31:0] r_run_copy10_j_281;
	reg  signed [31:0] r_run_copy0_j_282;
	reg  signed [31:0] r_run_copy1_j_283;
	reg  signed [31:0] r_run_copy2_j_284;
	reg  signed [31:0] r_run_copy3_j_285;
	reg  signed [31:0] r_run_copy4_j_286;
	reg  signed [31:0] r_run_copy5_j_287;
	reg  signed [31:0] r_run_copy6_j_288;
	reg  signed [31:0] r_run_copy7_j_289;
	reg  signed [31:0] r_run_copy8_j_290;
	reg  signed [31:0] r_run_copy9_j_291;
	reg  signed [31:0] r_run_copy10_j_292;
	reg  signed [31:0] r_run_copy0_j_293;
	reg  signed [31:0] r_run_copy1_j_294;
	reg  signed [31:0] r_run_copy2_j_295;
	reg  signed [31:0] r_run_copy3_j_296;
	reg  signed [31:0] r_run_copy4_j_297;
	reg  signed [31:0] r_run_copy5_j_298;
	reg  signed [31:0] r_run_copy6_j_299;
	reg  signed [31:0] r_run_copy7_j_300;
	reg  signed [31:0] r_run_copy8_j_301;
	reg  signed [31:0] r_run_copy9_j_302;
	reg  signed [31:0] r_run_copy10_j_303;
	reg  signed [31:0] r_run_copy0_j_304;
	reg  signed [31:0] r_run_copy0_j_305;
	reg  signed [31:0] r_run_copy1_j_306;
	reg  signed [31:0] r_run_copy0_j_307;
	reg  signed [31:0] r_run_copy1_j_308;
	reg  signed [31:0] r_run_copy0_j_309;
	reg  signed [31:0] r_run_copy1_j_310;
	reg  signed [31:0] r_run_copy0_j_311;
	reg  signed [31:0] r_run_copy1_j_312;
	reg  signed [31:0] r_run_copy0_j_313;
	reg  signed [31:0] r_run_copy1_j_314;
	reg  signed [31:0] r_run_copy0_j_315;
	reg  signed [31:0] r_run_copy1_j_316;
	reg  signed [31:0] r_run_copy0_j_317;
	reg  signed [31:0] r_run_copy1_j_318;
	reg  signed [31:0] r_run_copy0_j_319;
	reg  signed [31:0] r_run_copy0_j_320;
	reg  signed [31:0] r_run_copy1_j_321;
	reg  signed [31:0] r_run_copy0_j_322;
	reg  signed [31:0] r_run_copy1_j_323;
	reg  signed [31:0] r_run_copy0_j_324;
	reg  signed [31:0] r_run_copy1_j_325;
	reg  signed [31:0] r_run_copy0_j_326;
	reg  signed [31:0] r_run_copy1_j_327;
	reg  signed [31:0] r_run_copy0_j_328;
	reg  signed [31:0] r_run_copy1_j_329;
	reg  signed [31:0] r_run_copy0_j_330;
	reg  signed [31:0] r_run_copy1_j_331;
	reg  signed [31:0] r_run_copy0_j_332;
	reg  signed [31:0] r_run_copy1_j_333;
	reg  signed [31:0] r_run_copy0_j_334;
	reg  signed [31:0] r_run_copy0_j_335;
	reg  signed [31:0] r_run_copy1_j_336;
	reg  signed [31:0] r_run_copy0_j_337;
	reg  signed [31:0] r_run_copy1_j_338;
	reg  signed [31:0] r_run_copy0_j_339;
	reg  signed [31:0] r_run_copy1_j_340;
	reg  signed [31:0] r_run_copy0_j_341;
	reg  signed [31:0] r_run_copy1_j_342;
	reg  signed [31:0] r_run_copy0_j_343;
	reg  signed [31:0] r_run_copy1_j_344;
	reg  signed [31:0] r_run_copy0_j_345;
	reg  signed [31:0] r_run_copy1_j_346;
	reg  signed [31:0] r_run_copy0_j_347;
	reg  signed [31:0] r_run_copy1_j_348;
	reg  signed [31:0] r_run_copy0_j_349;
	reg  signed [31:0] r_run_copy0_j_350;
	reg  signed [31:0] r_run_copy1_j_351;
	reg  signed [31:0] r_run_copy0_j_352;
	reg  signed [31:0] r_run_copy1_j_353;
	reg  signed [31:0] r_run_copy0_j_354;
	reg  signed [31:0] r_run_copy1_j_355;
	reg  signed [31:0] r_run_copy0_j_356;
	reg  signed [31:0] r_run_copy1_j_357;
	reg  signed [31:0] r_run_copy0_j_358;
	reg  signed [31:0] r_run_copy1_j_359;
	reg  signed [31:0] r_run_copy0_j_360;
	reg  signed [31:0] r_run_copy1_j_361;
	reg  signed [31:0] r_run_copy0_j_362;
	reg  signed [31:0] r_run_copy1_j_363;
	reg                r_sub19_run_req;
	wire               w_sub19_run_busy;
	wire signed [14:0] w_sub19_T_addr;
	reg  signed [14:0] r_sub19_T_addr;
	wire        [31:0] w_sub19_T_datain;
	reg         [31:0] r_sub19_T_datain;
	wire        [31:0] w_sub19_T_dataout;
	wire               w_sub19_T_r_w;
	reg                r_sub19_T_r_w;
	wire signed [14:0] w_sub19_V_addr;
	reg  signed [14:0] r_sub19_V_addr;
	wire        [31:0] w_sub19_V_datain;
	reg         [31:0] r_sub19_V_datain;
	wire        [31:0] w_sub19_V_dataout;
	wire               w_sub19_V_r_w;
	reg                r_sub19_V_r_w;
	wire signed [14:0] w_sub19_U_addr;
	reg  signed [14:0] r_sub19_U_addr;
	wire        [31:0] w_sub19_U_datain;
	reg         [31:0] r_sub19_U_datain;
	wire        [31:0] w_sub19_U_dataout;
	wire               w_sub19_U_r_w;
	reg                r_sub19_U_r_w;
	wire signed [14:0] w_sub19_result_addr;
	reg  signed [14:0] r_sub19_result_addr;
	wire        [31:0] w_sub19_result_datain;
	reg         [31:0] r_sub19_result_datain;
	wire        [31:0] w_sub19_result_dataout;
	wire               w_sub19_result_r_w;
	reg                r_sub19_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [14:0] w_sub12_T_addr;
	reg  signed [14:0] r_sub12_T_addr;
	wire        [31:0] w_sub12_T_datain;
	reg         [31:0] r_sub12_T_datain;
	wire        [31:0] w_sub12_T_dataout;
	wire               w_sub12_T_r_w;
	reg                r_sub12_T_r_w;
	wire signed [14:0] w_sub12_V_addr;
	reg  signed [14:0] r_sub12_V_addr;
	wire        [31:0] w_sub12_V_datain;
	reg         [31:0] r_sub12_V_datain;
	wire        [31:0] w_sub12_V_dataout;
	wire               w_sub12_V_r_w;
	reg                r_sub12_V_r_w;
	wire signed [14:0] w_sub12_U_addr;
	reg  signed [14:0] r_sub12_U_addr;
	wire        [31:0] w_sub12_U_datain;
	reg         [31:0] r_sub12_U_datain;
	wire        [31:0] w_sub12_U_dataout;
	wire               w_sub12_U_r_w;
	reg                r_sub12_U_r_w;
	wire signed [14:0] w_sub12_result_addr;
	reg  signed [14:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [14:0] w_sub11_T_addr;
	reg  signed [14:0] r_sub11_T_addr;
	wire        [31:0] w_sub11_T_datain;
	reg         [31:0] r_sub11_T_datain;
	wire        [31:0] w_sub11_T_dataout;
	wire               w_sub11_T_r_w;
	reg                r_sub11_T_r_w;
	wire signed [14:0] w_sub11_V_addr;
	reg  signed [14:0] r_sub11_V_addr;
	wire        [31:0] w_sub11_V_datain;
	reg         [31:0] r_sub11_V_datain;
	wire        [31:0] w_sub11_V_dataout;
	wire               w_sub11_V_r_w;
	reg                r_sub11_V_r_w;
	wire signed [14:0] w_sub11_U_addr;
	reg  signed [14:0] r_sub11_U_addr;
	wire        [31:0] w_sub11_U_datain;
	reg         [31:0] r_sub11_U_datain;
	wire        [31:0] w_sub11_U_dataout;
	wire               w_sub11_U_r_w;
	reg                r_sub11_U_r_w;
	wire signed [14:0] w_sub11_result_addr;
	reg  signed [14:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [14:0] w_sub14_T_addr;
	reg  signed [14:0] r_sub14_T_addr;
	wire        [31:0] w_sub14_T_datain;
	reg         [31:0] r_sub14_T_datain;
	wire        [31:0] w_sub14_T_dataout;
	wire               w_sub14_T_r_w;
	reg                r_sub14_T_r_w;
	wire signed [14:0] w_sub14_V_addr;
	reg  signed [14:0] r_sub14_V_addr;
	wire        [31:0] w_sub14_V_datain;
	reg         [31:0] r_sub14_V_datain;
	wire        [31:0] w_sub14_V_dataout;
	wire               w_sub14_V_r_w;
	reg                r_sub14_V_r_w;
	wire signed [14:0] w_sub14_U_addr;
	reg  signed [14:0] r_sub14_U_addr;
	wire        [31:0] w_sub14_U_datain;
	reg         [31:0] r_sub14_U_datain;
	wire        [31:0] w_sub14_U_dataout;
	wire               w_sub14_U_r_w;
	reg                r_sub14_U_r_w;
	wire signed [14:0] w_sub14_result_addr;
	reg  signed [14:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [14:0] w_sub13_T_addr;
	reg  signed [14:0] r_sub13_T_addr;
	wire        [31:0] w_sub13_T_datain;
	reg         [31:0] r_sub13_T_datain;
	wire        [31:0] w_sub13_T_dataout;
	wire               w_sub13_T_r_w;
	reg                r_sub13_T_r_w;
	wire signed [14:0] w_sub13_V_addr;
	reg  signed [14:0] r_sub13_V_addr;
	wire        [31:0] w_sub13_V_datain;
	reg         [31:0] r_sub13_V_datain;
	wire        [31:0] w_sub13_V_dataout;
	wire               w_sub13_V_r_w;
	reg                r_sub13_V_r_w;
	wire signed [14:0] w_sub13_U_addr;
	reg  signed [14:0] r_sub13_U_addr;
	wire        [31:0] w_sub13_U_datain;
	reg         [31:0] r_sub13_U_datain;
	wire        [31:0] w_sub13_U_dataout;
	wire               w_sub13_U_r_w;
	reg                r_sub13_U_r_w;
	wire signed [14:0] w_sub13_result_addr;
	reg  signed [14:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub16_run_req;
	wire               w_sub16_run_busy;
	wire signed [14:0] w_sub16_T_addr;
	reg  signed [14:0] r_sub16_T_addr;
	wire        [31:0] w_sub16_T_datain;
	reg         [31:0] r_sub16_T_datain;
	wire        [31:0] w_sub16_T_dataout;
	wire               w_sub16_T_r_w;
	reg                r_sub16_T_r_w;
	wire signed [14:0] w_sub16_V_addr;
	reg  signed [14:0] r_sub16_V_addr;
	wire        [31:0] w_sub16_V_datain;
	reg         [31:0] r_sub16_V_datain;
	wire        [31:0] w_sub16_V_dataout;
	wire               w_sub16_V_r_w;
	reg                r_sub16_V_r_w;
	wire signed [14:0] w_sub16_U_addr;
	reg  signed [14:0] r_sub16_U_addr;
	wire        [31:0] w_sub16_U_datain;
	reg         [31:0] r_sub16_U_datain;
	wire        [31:0] w_sub16_U_dataout;
	wire               w_sub16_U_r_w;
	reg                r_sub16_U_r_w;
	wire signed [14:0] w_sub16_result_addr;
	reg  signed [14:0] r_sub16_result_addr;
	wire        [31:0] w_sub16_result_datain;
	reg         [31:0] r_sub16_result_datain;
	wire        [31:0] w_sub16_result_dataout;
	wire               w_sub16_result_r_w;
	reg                r_sub16_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [14:0] w_sub15_T_addr;
	reg  signed [14:0] r_sub15_T_addr;
	wire        [31:0] w_sub15_T_datain;
	reg         [31:0] r_sub15_T_datain;
	wire        [31:0] w_sub15_T_dataout;
	wire               w_sub15_T_r_w;
	reg                r_sub15_T_r_w;
	wire signed [14:0] w_sub15_V_addr;
	reg  signed [14:0] r_sub15_V_addr;
	wire        [31:0] w_sub15_V_datain;
	reg         [31:0] r_sub15_V_datain;
	wire        [31:0] w_sub15_V_dataout;
	wire               w_sub15_V_r_w;
	reg                r_sub15_V_r_w;
	wire signed [14:0] w_sub15_U_addr;
	reg  signed [14:0] r_sub15_U_addr;
	wire        [31:0] w_sub15_U_datain;
	reg         [31:0] r_sub15_U_datain;
	wire        [31:0] w_sub15_U_dataout;
	wire               w_sub15_U_r_w;
	reg                r_sub15_U_r_w;
	wire signed [14:0] w_sub15_result_addr;
	reg  signed [14:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub18_run_req;
	wire               w_sub18_run_busy;
	wire signed [14:0] w_sub18_T_addr;
	reg  signed [14:0] r_sub18_T_addr;
	wire        [31:0] w_sub18_T_datain;
	reg         [31:0] r_sub18_T_datain;
	wire        [31:0] w_sub18_T_dataout;
	wire               w_sub18_T_r_w;
	reg                r_sub18_T_r_w;
	wire signed [14:0] w_sub18_V_addr;
	reg  signed [14:0] r_sub18_V_addr;
	wire        [31:0] w_sub18_V_datain;
	reg         [31:0] r_sub18_V_datain;
	wire        [31:0] w_sub18_V_dataout;
	wire               w_sub18_V_r_w;
	reg                r_sub18_V_r_w;
	wire signed [14:0] w_sub18_U_addr;
	reg  signed [14:0] r_sub18_U_addr;
	wire        [31:0] w_sub18_U_datain;
	reg         [31:0] r_sub18_U_datain;
	wire        [31:0] w_sub18_U_dataout;
	wire               w_sub18_U_r_w;
	reg                r_sub18_U_r_w;
	wire signed [14:0] w_sub18_result_addr;
	reg  signed [14:0] r_sub18_result_addr;
	wire        [31:0] w_sub18_result_datain;
	reg         [31:0] r_sub18_result_datain;
	wire        [31:0] w_sub18_result_dataout;
	wire               w_sub18_result_r_w;
	reg                r_sub18_result_r_w;
	reg                r_sub17_run_req;
	wire               w_sub17_run_busy;
	wire signed [14:0] w_sub17_T_addr;
	reg  signed [14:0] r_sub17_T_addr;
	wire        [31:0] w_sub17_T_datain;
	reg         [31:0] r_sub17_T_datain;
	wire        [31:0] w_sub17_T_dataout;
	wire               w_sub17_T_r_w;
	reg                r_sub17_T_r_w;
	wire signed [14:0] w_sub17_V_addr;
	reg  signed [14:0] r_sub17_V_addr;
	wire        [31:0] w_sub17_V_datain;
	reg         [31:0] r_sub17_V_datain;
	wire        [31:0] w_sub17_V_dataout;
	wire               w_sub17_V_r_w;
	reg                r_sub17_V_r_w;
	wire signed [14:0] w_sub17_U_addr;
	reg  signed [14:0] r_sub17_U_addr;
	wire        [31:0] w_sub17_U_datain;
	reg         [31:0] r_sub17_U_datain;
	wire        [31:0] w_sub17_U_dataout;
	wire               w_sub17_U_r_w;
	reg                r_sub17_U_r_w;
	wire signed [14:0] w_sub17_result_addr;
	reg  signed [14:0] r_sub17_result_addr;
	wire        [31:0] w_sub17_result_datain;
	reg         [31:0] r_sub17_result_datain;
	wire        [31:0] w_sub17_result_dataout;
	wire               w_sub17_result_r_w;
	reg                r_sub17_result_r_w;
	reg                r_sub20_run_req;
	wire               w_sub20_run_busy;
	wire signed [14:0] w_sub20_T_addr;
	reg  signed [14:0] r_sub20_T_addr;
	wire        [31:0] w_sub20_T_datain;
	reg         [31:0] r_sub20_T_datain;
	wire        [31:0] w_sub20_T_dataout;
	wire               w_sub20_T_r_w;
	reg                r_sub20_T_r_w;
	wire signed [14:0] w_sub20_V_addr;
	reg  signed [14:0] r_sub20_V_addr;
	wire        [31:0] w_sub20_V_datain;
	reg         [31:0] r_sub20_V_datain;
	wire        [31:0] w_sub20_V_dataout;
	wire               w_sub20_V_r_w;
	reg                r_sub20_V_r_w;
	wire signed [14:0] w_sub20_U_addr;
	reg  signed [14:0] r_sub20_U_addr;
	wire        [31:0] w_sub20_U_datain;
	reg         [31:0] r_sub20_U_datain;
	wire        [31:0] w_sub20_U_dataout;
	wire               w_sub20_U_r_w;
	reg                r_sub20_U_r_w;
	wire signed [14:0] w_sub20_result_addr;
	reg  signed [14:0] r_sub20_result_addr;
	wire        [31:0] w_sub20_result_datain;
	reg         [31:0] r_sub20_result_datain;
	wire        [31:0] w_sub20_result_dataout;
	wire               w_sub20_result_r_w;
	reg                r_sub20_result_r_w;
	reg                r_sub21_run_req;
	wire               w_sub21_run_busy;
	wire signed [14:0] w_sub21_T_addr;
	reg  signed [14:0] r_sub21_T_addr;
	wire        [31:0] w_sub21_T_datain;
	reg         [31:0] r_sub21_T_datain;
	wire        [31:0] w_sub21_T_dataout;
	wire               w_sub21_T_r_w;
	reg                r_sub21_T_r_w;
	wire signed [14:0] w_sub21_V_addr;
	reg  signed [14:0] r_sub21_V_addr;
	wire        [31:0] w_sub21_V_datain;
	reg         [31:0] r_sub21_V_datain;
	wire        [31:0] w_sub21_V_dataout;
	wire               w_sub21_V_r_w;
	reg                r_sub21_V_r_w;
	wire signed [14:0] w_sub21_U_addr;
	reg  signed [14:0] r_sub21_U_addr;
	wire        [31:0] w_sub21_U_datain;
	reg         [31:0] r_sub21_U_datain;
	wire        [31:0] w_sub21_U_dataout;
	wire               w_sub21_U_r_w;
	reg                r_sub21_U_r_w;
	wire signed [14:0] w_sub21_result_addr;
	reg  signed [14:0] r_sub21_result_addr;
	wire        [31:0] w_sub21_result_datain;
	reg         [31:0] r_sub21_result_datain;
	wire        [31:0] w_sub21_result_dataout;
	wire               w_sub21_result_r_w;
	reg                r_sub21_result_r_w;
	reg                r_sub28_run_req;
	wire               w_sub28_run_busy;
	wire signed [14:0] w_sub28_T_addr;
	reg  signed [14:0] r_sub28_T_addr;
	wire        [31:0] w_sub28_T_datain;
	reg         [31:0] r_sub28_T_datain;
	wire        [31:0] w_sub28_T_dataout;
	wire               w_sub28_T_r_w;
	reg                r_sub28_T_r_w;
	wire signed [14:0] w_sub28_V_addr;
	reg  signed [14:0] r_sub28_V_addr;
	wire        [31:0] w_sub28_V_datain;
	reg         [31:0] r_sub28_V_datain;
	wire        [31:0] w_sub28_V_dataout;
	wire               w_sub28_V_r_w;
	reg                r_sub28_V_r_w;
	wire signed [14:0] w_sub28_U_addr;
	reg  signed [14:0] r_sub28_U_addr;
	wire        [31:0] w_sub28_U_datain;
	reg         [31:0] r_sub28_U_datain;
	wire        [31:0] w_sub28_U_dataout;
	wire               w_sub28_U_r_w;
	reg                r_sub28_U_r_w;
	wire signed [14:0] w_sub28_result_addr;
	reg  signed [14:0] r_sub28_result_addr;
	wire        [31:0] w_sub28_result_datain;
	reg         [31:0] r_sub28_result_datain;
	wire        [31:0] w_sub28_result_dataout;
	wire               w_sub28_result_r_w;
	reg                r_sub28_result_r_w;
	reg                r_sub29_run_req;
	wire               w_sub29_run_busy;
	wire signed [14:0] w_sub29_T_addr;
	reg  signed [14:0] r_sub29_T_addr;
	wire        [31:0] w_sub29_T_datain;
	reg         [31:0] r_sub29_T_datain;
	wire        [31:0] w_sub29_T_dataout;
	wire               w_sub29_T_r_w;
	reg                r_sub29_T_r_w;
	wire signed [14:0] w_sub29_V_addr;
	reg  signed [14:0] r_sub29_V_addr;
	wire        [31:0] w_sub29_V_datain;
	reg         [31:0] r_sub29_V_datain;
	wire        [31:0] w_sub29_V_dataout;
	wire               w_sub29_V_r_w;
	reg                r_sub29_V_r_w;
	wire signed [14:0] w_sub29_U_addr;
	reg  signed [14:0] r_sub29_U_addr;
	wire        [31:0] w_sub29_U_datain;
	reg         [31:0] r_sub29_U_datain;
	wire        [31:0] w_sub29_U_dataout;
	wire               w_sub29_U_r_w;
	reg                r_sub29_U_r_w;
	wire signed [14:0] w_sub29_result_addr;
	reg  signed [14:0] r_sub29_result_addr;
	wire        [31:0] w_sub29_result_datain;
	reg         [31:0] r_sub29_result_datain;
	wire        [31:0] w_sub29_result_dataout;
	wire               w_sub29_result_r_w;
	reg                r_sub29_result_r_w;
	reg                r_sub26_run_req;
	wire               w_sub26_run_busy;
	wire signed [14:0] w_sub26_T_addr;
	reg  signed [14:0] r_sub26_T_addr;
	wire        [31:0] w_sub26_T_datain;
	reg         [31:0] r_sub26_T_datain;
	wire        [31:0] w_sub26_T_dataout;
	wire               w_sub26_T_r_w;
	reg                r_sub26_T_r_w;
	wire signed [14:0] w_sub26_V_addr;
	reg  signed [14:0] r_sub26_V_addr;
	wire        [31:0] w_sub26_V_datain;
	reg         [31:0] r_sub26_V_datain;
	wire        [31:0] w_sub26_V_dataout;
	wire               w_sub26_V_r_w;
	reg                r_sub26_V_r_w;
	wire signed [14:0] w_sub26_U_addr;
	reg  signed [14:0] r_sub26_U_addr;
	wire        [31:0] w_sub26_U_datain;
	reg         [31:0] r_sub26_U_datain;
	wire        [31:0] w_sub26_U_dataout;
	wire               w_sub26_U_r_w;
	reg                r_sub26_U_r_w;
	wire signed [14:0] w_sub26_result_addr;
	reg  signed [14:0] r_sub26_result_addr;
	wire        [31:0] w_sub26_result_datain;
	reg         [31:0] r_sub26_result_datain;
	wire        [31:0] w_sub26_result_dataout;
	wire               w_sub26_result_r_w;
	reg                r_sub26_result_r_w;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [14:0] w_sub09_T_addr;
	reg  signed [14:0] r_sub09_T_addr;
	wire        [31:0] w_sub09_T_datain;
	reg         [31:0] r_sub09_T_datain;
	wire        [31:0] w_sub09_T_dataout;
	wire               w_sub09_T_r_w;
	reg                r_sub09_T_r_w;
	wire signed [14:0] w_sub09_V_addr;
	reg  signed [14:0] r_sub09_V_addr;
	wire        [31:0] w_sub09_V_datain;
	reg         [31:0] r_sub09_V_datain;
	wire        [31:0] w_sub09_V_dataout;
	wire               w_sub09_V_r_w;
	reg                r_sub09_V_r_w;
	wire signed [14:0] w_sub09_U_addr;
	reg  signed [14:0] r_sub09_U_addr;
	wire        [31:0] w_sub09_U_datain;
	reg         [31:0] r_sub09_U_datain;
	wire        [31:0] w_sub09_U_dataout;
	wire               w_sub09_U_r_w;
	reg                r_sub09_U_r_w;
	wire signed [14:0] w_sub09_result_addr;
	reg  signed [14:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub27_run_req;
	wire               w_sub27_run_busy;
	wire signed [14:0] w_sub27_T_addr;
	reg  signed [14:0] r_sub27_T_addr;
	wire        [31:0] w_sub27_T_datain;
	reg         [31:0] r_sub27_T_datain;
	wire        [31:0] w_sub27_T_dataout;
	wire               w_sub27_T_r_w;
	reg                r_sub27_T_r_w;
	wire signed [14:0] w_sub27_V_addr;
	reg  signed [14:0] r_sub27_V_addr;
	wire        [31:0] w_sub27_V_datain;
	reg         [31:0] r_sub27_V_datain;
	wire        [31:0] w_sub27_V_dataout;
	wire               w_sub27_V_r_w;
	reg                r_sub27_V_r_w;
	wire signed [14:0] w_sub27_U_addr;
	reg  signed [14:0] r_sub27_U_addr;
	wire        [31:0] w_sub27_U_datain;
	reg         [31:0] r_sub27_U_datain;
	wire        [31:0] w_sub27_U_dataout;
	wire               w_sub27_U_r_w;
	reg                r_sub27_U_r_w;
	wire signed [14:0] w_sub27_result_addr;
	reg  signed [14:0] r_sub27_result_addr;
	wire        [31:0] w_sub27_result_datain;
	reg         [31:0] r_sub27_result_datain;
	wire        [31:0] w_sub27_result_dataout;
	wire               w_sub27_result_r_w;
	reg                r_sub27_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [14:0] w_sub08_T_addr;
	reg  signed [14:0] r_sub08_T_addr;
	wire        [31:0] w_sub08_T_datain;
	reg         [31:0] r_sub08_T_datain;
	wire        [31:0] w_sub08_T_dataout;
	wire               w_sub08_T_r_w;
	reg                r_sub08_T_r_w;
	wire signed [14:0] w_sub08_V_addr;
	reg  signed [14:0] r_sub08_V_addr;
	wire        [31:0] w_sub08_V_datain;
	reg         [31:0] r_sub08_V_datain;
	wire        [31:0] w_sub08_V_dataout;
	wire               w_sub08_V_r_w;
	reg                r_sub08_V_r_w;
	wire signed [14:0] w_sub08_U_addr;
	reg  signed [14:0] r_sub08_U_addr;
	wire        [31:0] w_sub08_U_datain;
	reg         [31:0] r_sub08_U_datain;
	wire        [31:0] w_sub08_U_dataout;
	wire               w_sub08_U_r_w;
	reg                r_sub08_U_r_w;
	wire signed [14:0] w_sub08_result_addr;
	reg  signed [14:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub24_run_req;
	wire               w_sub24_run_busy;
	wire signed [14:0] w_sub24_T_addr;
	reg  signed [14:0] r_sub24_T_addr;
	wire        [31:0] w_sub24_T_datain;
	reg         [31:0] r_sub24_T_datain;
	wire        [31:0] w_sub24_T_dataout;
	wire               w_sub24_T_r_w;
	reg                r_sub24_T_r_w;
	wire signed [14:0] w_sub24_V_addr;
	reg  signed [14:0] r_sub24_V_addr;
	wire        [31:0] w_sub24_V_datain;
	reg         [31:0] r_sub24_V_datain;
	wire        [31:0] w_sub24_V_dataout;
	wire               w_sub24_V_r_w;
	reg                r_sub24_V_r_w;
	wire signed [14:0] w_sub24_U_addr;
	reg  signed [14:0] r_sub24_U_addr;
	wire        [31:0] w_sub24_U_datain;
	reg         [31:0] r_sub24_U_datain;
	wire        [31:0] w_sub24_U_dataout;
	wire               w_sub24_U_r_w;
	reg                r_sub24_U_r_w;
	wire signed [14:0] w_sub24_result_addr;
	reg  signed [14:0] r_sub24_result_addr;
	wire        [31:0] w_sub24_result_datain;
	reg         [31:0] r_sub24_result_datain;
	wire        [31:0] w_sub24_result_dataout;
	wire               w_sub24_result_r_w;
	reg                r_sub24_result_r_w;
	reg                r_sub25_run_req;
	wire               w_sub25_run_busy;
	wire signed [14:0] w_sub25_T_addr;
	reg  signed [14:0] r_sub25_T_addr;
	wire        [31:0] w_sub25_T_datain;
	reg         [31:0] r_sub25_T_datain;
	wire        [31:0] w_sub25_T_dataout;
	wire               w_sub25_T_r_w;
	reg                r_sub25_T_r_w;
	wire signed [14:0] w_sub25_V_addr;
	reg  signed [14:0] r_sub25_V_addr;
	wire        [31:0] w_sub25_V_datain;
	reg         [31:0] r_sub25_V_datain;
	wire        [31:0] w_sub25_V_dataout;
	wire               w_sub25_V_r_w;
	reg                r_sub25_V_r_w;
	wire signed [14:0] w_sub25_U_addr;
	reg  signed [14:0] r_sub25_U_addr;
	wire        [31:0] w_sub25_U_datain;
	reg         [31:0] r_sub25_U_datain;
	wire        [31:0] w_sub25_U_dataout;
	wire               w_sub25_U_r_w;
	reg                r_sub25_U_r_w;
	wire signed [14:0] w_sub25_result_addr;
	reg  signed [14:0] r_sub25_result_addr;
	wire        [31:0] w_sub25_result_datain;
	reg         [31:0] r_sub25_result_datain;
	wire        [31:0] w_sub25_result_dataout;
	wire               w_sub25_result_r_w;
	reg                r_sub25_result_r_w;
	reg                r_sub22_run_req;
	wire               w_sub22_run_busy;
	wire signed [14:0] w_sub22_T_addr;
	reg  signed [14:0] r_sub22_T_addr;
	wire        [31:0] w_sub22_T_datain;
	reg         [31:0] r_sub22_T_datain;
	wire        [31:0] w_sub22_T_dataout;
	wire               w_sub22_T_r_w;
	reg                r_sub22_T_r_w;
	wire signed [14:0] w_sub22_V_addr;
	reg  signed [14:0] r_sub22_V_addr;
	wire        [31:0] w_sub22_V_datain;
	reg         [31:0] r_sub22_V_datain;
	wire        [31:0] w_sub22_V_dataout;
	wire               w_sub22_V_r_w;
	reg                r_sub22_V_r_w;
	wire signed [14:0] w_sub22_U_addr;
	reg  signed [14:0] r_sub22_U_addr;
	wire        [31:0] w_sub22_U_datain;
	reg         [31:0] r_sub22_U_datain;
	wire        [31:0] w_sub22_U_dataout;
	wire               w_sub22_U_r_w;
	reg                r_sub22_U_r_w;
	wire signed [14:0] w_sub22_result_addr;
	reg  signed [14:0] r_sub22_result_addr;
	wire        [31:0] w_sub22_result_datain;
	reg         [31:0] r_sub22_result_datain;
	wire        [31:0] w_sub22_result_dataout;
	wire               w_sub22_result_r_w;
	reg                r_sub22_result_r_w;
	reg                r_sub23_run_req;
	wire               w_sub23_run_busy;
	wire signed [14:0] w_sub23_T_addr;
	reg  signed [14:0] r_sub23_T_addr;
	wire        [31:0] w_sub23_T_datain;
	reg         [31:0] r_sub23_T_datain;
	wire        [31:0] w_sub23_T_dataout;
	wire               w_sub23_T_r_w;
	reg                r_sub23_T_r_w;
	wire signed [14:0] w_sub23_V_addr;
	reg  signed [14:0] r_sub23_V_addr;
	wire        [31:0] w_sub23_V_datain;
	reg         [31:0] r_sub23_V_datain;
	wire        [31:0] w_sub23_V_dataout;
	wire               w_sub23_V_r_w;
	reg                r_sub23_V_r_w;
	wire signed [14:0] w_sub23_U_addr;
	reg  signed [14:0] r_sub23_U_addr;
	wire        [31:0] w_sub23_U_datain;
	reg         [31:0] r_sub23_U_datain;
	wire        [31:0] w_sub23_U_dataout;
	wire               w_sub23_U_r_w;
	reg                r_sub23_U_r_w;
	wire signed [14:0] w_sub23_result_addr;
	reg  signed [14:0] r_sub23_result_addr;
	wire        [31:0] w_sub23_result_datain;
	reg         [31:0] r_sub23_result_datain;
	wire        [31:0] w_sub23_result_dataout;
	wire               w_sub23_result_r_w;
	reg                r_sub23_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [14:0] w_sub03_T_addr;
	reg  signed [14:0] r_sub03_T_addr;
	wire        [31:0] w_sub03_T_datain;
	reg         [31:0] r_sub03_T_datain;
	wire        [31:0] w_sub03_T_dataout;
	wire               w_sub03_T_r_w;
	reg                r_sub03_T_r_w;
	wire signed [14:0] w_sub03_V_addr;
	reg  signed [14:0] r_sub03_V_addr;
	wire        [31:0] w_sub03_V_datain;
	reg         [31:0] r_sub03_V_datain;
	wire        [31:0] w_sub03_V_dataout;
	wire               w_sub03_V_r_w;
	reg                r_sub03_V_r_w;
	wire signed [14:0] w_sub03_U_addr;
	reg  signed [14:0] r_sub03_U_addr;
	wire        [31:0] w_sub03_U_datain;
	reg         [31:0] r_sub03_U_datain;
	wire        [31:0] w_sub03_U_dataout;
	wire               w_sub03_U_r_w;
	reg                r_sub03_U_r_w;
	wire signed [14:0] w_sub03_result_addr;
	reg  signed [14:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [14:0] w_sub02_T_addr;
	reg  signed [14:0] r_sub02_T_addr;
	wire        [31:0] w_sub02_T_datain;
	reg         [31:0] r_sub02_T_datain;
	wire        [31:0] w_sub02_T_dataout;
	wire               w_sub02_T_r_w;
	reg                r_sub02_T_r_w;
	wire signed [14:0] w_sub02_V_addr;
	reg  signed [14:0] r_sub02_V_addr;
	wire        [31:0] w_sub02_V_datain;
	reg         [31:0] r_sub02_V_datain;
	wire        [31:0] w_sub02_V_dataout;
	wire               w_sub02_V_r_w;
	reg                r_sub02_V_r_w;
	wire signed [14:0] w_sub02_U_addr;
	reg  signed [14:0] r_sub02_U_addr;
	wire        [31:0] w_sub02_U_datain;
	reg         [31:0] r_sub02_U_datain;
	wire        [31:0] w_sub02_U_dataout;
	wire               w_sub02_U_r_w;
	reg                r_sub02_U_r_w;
	wire signed [14:0] w_sub02_result_addr;
	reg  signed [14:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [14:0] w_sub01_T_addr;
	reg  signed [14:0] r_sub01_T_addr;
	wire        [31:0] w_sub01_T_datain;
	reg         [31:0] r_sub01_T_datain;
	wire        [31:0] w_sub01_T_dataout;
	wire               w_sub01_T_r_w;
	reg                r_sub01_T_r_w;
	wire signed [14:0] w_sub01_V_addr;
	reg  signed [14:0] r_sub01_V_addr;
	wire        [31:0] w_sub01_V_datain;
	reg         [31:0] r_sub01_V_datain;
	wire        [31:0] w_sub01_V_dataout;
	wire               w_sub01_V_r_w;
	reg                r_sub01_V_r_w;
	wire signed [14:0] w_sub01_U_addr;
	reg  signed [14:0] r_sub01_U_addr;
	wire        [31:0] w_sub01_U_datain;
	reg         [31:0] r_sub01_U_datain;
	wire        [31:0] w_sub01_U_dataout;
	wire               w_sub01_U_r_w;
	reg                r_sub01_U_r_w;
	wire signed [14:0] w_sub01_result_addr;
	reg  signed [14:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [14:0] w_sub00_T_addr;
	reg  signed [14:0] r_sub00_T_addr;
	wire        [31:0] w_sub00_T_datain;
	reg         [31:0] r_sub00_T_datain;
	wire        [31:0] w_sub00_T_dataout;
	wire               w_sub00_T_r_w;
	reg                r_sub00_T_r_w;
	wire signed [14:0] w_sub00_V_addr;
	reg  signed [14:0] r_sub00_V_addr;
	wire        [31:0] w_sub00_V_datain;
	reg         [31:0] r_sub00_V_datain;
	wire        [31:0] w_sub00_V_dataout;
	wire               w_sub00_V_r_w;
	reg                r_sub00_V_r_w;
	wire signed [14:0] w_sub00_U_addr;
	reg  signed [14:0] r_sub00_U_addr;
	wire        [31:0] w_sub00_U_datain;
	reg         [31:0] r_sub00_U_datain;
	wire        [31:0] w_sub00_U_dataout;
	wire               w_sub00_U_r_w;
	reg                r_sub00_U_r_w;
	wire signed [14:0] w_sub00_result_addr;
	reg  signed [14:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [14:0] w_sub07_T_addr;
	reg  signed [14:0] r_sub07_T_addr;
	wire        [31:0] w_sub07_T_datain;
	reg         [31:0] r_sub07_T_datain;
	wire        [31:0] w_sub07_T_dataout;
	wire               w_sub07_T_r_w;
	reg                r_sub07_T_r_w;
	wire signed [14:0] w_sub07_V_addr;
	reg  signed [14:0] r_sub07_V_addr;
	wire        [31:0] w_sub07_V_datain;
	reg         [31:0] r_sub07_V_datain;
	wire        [31:0] w_sub07_V_dataout;
	wire               w_sub07_V_r_w;
	reg                r_sub07_V_r_w;
	wire signed [14:0] w_sub07_U_addr;
	reg  signed [14:0] r_sub07_U_addr;
	wire        [31:0] w_sub07_U_datain;
	reg         [31:0] r_sub07_U_datain;
	wire        [31:0] w_sub07_U_dataout;
	wire               w_sub07_U_r_w;
	reg                r_sub07_U_r_w;
	wire signed [14:0] w_sub07_result_addr;
	reg  signed [14:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [14:0] w_sub06_T_addr;
	reg  signed [14:0] r_sub06_T_addr;
	wire        [31:0] w_sub06_T_datain;
	reg         [31:0] r_sub06_T_datain;
	wire        [31:0] w_sub06_T_dataout;
	wire               w_sub06_T_r_w;
	reg                r_sub06_T_r_w;
	wire signed [14:0] w_sub06_V_addr;
	reg  signed [14:0] r_sub06_V_addr;
	wire        [31:0] w_sub06_V_datain;
	reg         [31:0] r_sub06_V_datain;
	wire        [31:0] w_sub06_V_dataout;
	wire               w_sub06_V_r_w;
	reg                r_sub06_V_r_w;
	wire signed [14:0] w_sub06_U_addr;
	reg  signed [14:0] r_sub06_U_addr;
	wire        [31:0] w_sub06_U_datain;
	reg         [31:0] r_sub06_U_datain;
	wire        [31:0] w_sub06_U_dataout;
	wire               w_sub06_U_r_w;
	reg                r_sub06_U_r_w;
	wire signed [14:0] w_sub06_result_addr;
	reg  signed [14:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [14:0] w_sub05_T_addr;
	reg  signed [14:0] r_sub05_T_addr;
	wire        [31:0] w_sub05_T_datain;
	reg         [31:0] r_sub05_T_datain;
	wire        [31:0] w_sub05_T_dataout;
	wire               w_sub05_T_r_w;
	reg                r_sub05_T_r_w;
	wire signed [14:0] w_sub05_V_addr;
	reg  signed [14:0] r_sub05_V_addr;
	wire        [31:0] w_sub05_V_datain;
	reg         [31:0] r_sub05_V_datain;
	wire        [31:0] w_sub05_V_dataout;
	wire               w_sub05_V_r_w;
	reg                r_sub05_V_r_w;
	wire signed [14:0] w_sub05_U_addr;
	reg  signed [14:0] r_sub05_U_addr;
	wire        [31:0] w_sub05_U_datain;
	reg         [31:0] r_sub05_U_datain;
	wire        [31:0] w_sub05_U_dataout;
	wire               w_sub05_U_r_w;
	reg                r_sub05_U_r_w;
	wire signed [14:0] w_sub05_result_addr;
	reg  signed [14:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [14:0] w_sub04_T_addr;
	reg  signed [14:0] r_sub04_T_addr;
	wire        [31:0] w_sub04_T_datain;
	reg         [31:0] r_sub04_T_datain;
	wire        [31:0] w_sub04_T_dataout;
	wire               w_sub04_T_r_w;
	reg                r_sub04_T_r_w;
	wire signed [14:0] w_sub04_V_addr;
	reg  signed [14:0] r_sub04_V_addr;
	wire        [31:0] w_sub04_V_datain;
	reg         [31:0] r_sub04_V_datain;
	wire        [31:0] w_sub04_V_dataout;
	wire               w_sub04_V_r_w;
	reg                r_sub04_V_r_w;
	wire signed [14:0] w_sub04_U_addr;
	reg  signed [14:0] r_sub04_U_addr;
	wire        [31:0] w_sub04_U_datain;
	reg         [31:0] r_sub04_U_datain;
	wire        [31:0] w_sub04_U_dataout;
	wire               w_sub04_U_r_w;
	reg                r_sub04_U_r_w;
	wire signed [14:0] w_sub04_result_addr;
	reg  signed [14:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [14:0] w_sub10_T_addr;
	reg  signed [14:0] r_sub10_T_addr;
	wire        [31:0] w_sub10_T_datain;
	reg         [31:0] r_sub10_T_datain;
	wire        [31:0] w_sub10_T_dataout;
	wire               w_sub10_T_r_w;
	reg                r_sub10_T_r_w;
	wire signed [14:0] w_sub10_V_addr;
	reg  signed [14:0] r_sub10_V_addr;
	wire        [31:0] w_sub10_V_datain;
	reg         [31:0] r_sub10_V_datain;
	wire        [31:0] w_sub10_V_dataout;
	wire               w_sub10_V_r_w;
	reg                r_sub10_V_r_w;
	wire signed [14:0] w_sub10_U_addr;
	reg  signed [14:0] r_sub10_U_addr;
	wire        [31:0] w_sub10_U_datain;
	reg         [31:0] r_sub10_U_datain;
	wire        [31:0] w_sub10_U_dataout;
	wire               w_sub10_U_r_w;
	reg                r_sub10_U_r_w;
	wire signed [14:0] w_sub10_result_addr;
	reg  signed [14:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg                r_sub31_run_req;
	wire               w_sub31_run_busy;
	wire signed [14:0] w_sub31_T_addr;
	reg  signed [14:0] r_sub31_T_addr;
	wire        [31:0] w_sub31_T_datain;
	reg         [31:0] r_sub31_T_datain;
	wire        [31:0] w_sub31_T_dataout;
	wire               w_sub31_T_r_w;
	reg                r_sub31_T_r_w;
	wire signed [14:0] w_sub31_V_addr;
	reg  signed [14:0] r_sub31_V_addr;
	wire        [31:0] w_sub31_V_datain;
	reg         [31:0] r_sub31_V_datain;
	wire        [31:0] w_sub31_V_dataout;
	wire               w_sub31_V_r_w;
	reg                r_sub31_V_r_w;
	wire signed [14:0] w_sub31_U_addr;
	reg  signed [14:0] r_sub31_U_addr;
	wire        [31:0] w_sub31_U_datain;
	reg         [31:0] r_sub31_U_datain;
	wire        [31:0] w_sub31_U_dataout;
	wire               w_sub31_U_r_w;
	reg                r_sub31_U_r_w;
	wire signed [14:0] w_sub31_result_addr;
	reg  signed [14:0] r_sub31_result_addr;
	wire        [31:0] w_sub31_result_datain;
	reg         [31:0] r_sub31_result_datain;
	wire        [31:0] w_sub31_result_dataout;
	wire               w_sub31_result_r_w;
	reg                r_sub31_result_r_w;
	reg                r_sub30_run_req;
	wire               w_sub30_run_busy;
	wire signed [14:0] w_sub30_T_addr;
	reg  signed [14:0] r_sub30_T_addr;
	wire        [31:0] w_sub30_T_datain;
	reg         [31:0] r_sub30_T_datain;
	wire        [31:0] w_sub30_T_dataout;
	wire               w_sub30_T_r_w;
	reg                r_sub30_T_r_w;
	wire signed [14:0] w_sub30_V_addr;
	reg  signed [14:0] r_sub30_V_addr;
	wire        [31:0] w_sub30_V_datain;
	reg         [31:0] r_sub30_V_datain;
	wire        [31:0] w_sub30_V_dataout;
	wire               w_sub30_V_r_w;
	reg                r_sub30_V_r_w;
	wire signed [14:0] w_sub30_U_addr;
	reg  signed [14:0] r_sub30_U_addr;
	wire        [31:0] w_sub30_U_datain;
	reg         [31:0] r_sub30_U_datain;
	wire        [31:0] w_sub30_U_dataout;
	wire               w_sub30_U_r_w;
	reg                r_sub30_U_r_w;
	wire signed [14:0] w_sub30_result_addr;
	reg  signed [14:0] r_sub30_result_addr;
	wire        [31:0] w_sub30_result_datain;
	reg         [31:0] r_sub30_result_datain;
	wire        [31:0] w_sub30_result_dataout;
	wire               w_sub30_result_r_w;
	reg                r_sub30_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire               w_sys_tmp12;
	wire               w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp15;
	wire               w_sys_tmp16;
	wire        [31:0] w_sys_tmp18;
	wire        [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire        [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp27;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp32;
	wire signed [31:0] w_sys_tmp33;
	wire        [31:0] w_sys_tmp36;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp45;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire        [31:0] w_sys_tmp128;
	wire               w_sys_tmp226;
	wire               w_sys_tmp227;
	wire signed [31:0] w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire               w_sys_tmp230;
	wire               w_sys_tmp231;
	wire signed [31:0] w_sys_tmp232;
	wire signed [31:0] w_sys_tmp235;
	wire signed [31:0] w_sys_tmp236;
	wire signed [31:0] w_sys_tmp237;
	wire        [31:0] w_sys_tmp238;
	wire signed [31:0] w_sys_tmp239;
	wire signed [31:0] w_sys_tmp240;
	wire signed [31:0] w_sys_tmp243;
	wire signed [31:0] w_sys_tmp244;
	wire        [31:0] w_sys_tmp246;
	wire signed [31:0] w_sys_tmp247;
	wire signed [31:0] w_sys_tmp248;
	wire signed [31:0] w_sys_tmp251;
	wire signed [31:0] w_sys_tmp252;
	wire        [31:0] w_sys_tmp254;
	wire signed [31:0] w_sys_tmp255;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp258;
	wire signed [31:0] w_sys_tmp259;
	wire signed [31:0] w_sys_tmp260;
	wire signed [31:0] w_sys_tmp261;
	wire signed [31:0] w_sys_tmp262;
	wire signed [31:0] w_sys_tmp263;
	wire signed [31:0] w_sys_tmp444;
	wire               w_sys_tmp445;
	wire               w_sys_tmp446;
	wire signed [31:0] w_sys_tmp447;
	wire signed [31:0] w_sys_tmp450;
	wire signed [31:0] w_sys_tmp451;
	wire signed [31:0] w_sys_tmp452;
	wire        [31:0] w_sys_tmp453;
	wire signed [31:0] w_sys_tmp454;
	wire signed [31:0] w_sys_tmp455;
	wire signed [31:0] w_sys_tmp458;
	wire signed [31:0] w_sys_tmp459;
	wire        [31:0] w_sys_tmp461;
	wire signed [31:0] w_sys_tmp462;
	wire signed [31:0] w_sys_tmp463;
	wire signed [31:0] w_sys_tmp466;
	wire signed [31:0] w_sys_tmp467;
	wire        [31:0] w_sys_tmp469;
	wire signed [31:0] w_sys_tmp470;
	wire signed [31:0] w_sys_tmp471;
	wire signed [31:0] w_sys_tmp473;
	wire signed [31:0] w_sys_tmp474;
	wire signed [31:0] w_sys_tmp475;
	wire signed [31:0] w_sys_tmp476;
	wire signed [31:0] w_sys_tmp477;
	wire signed [31:0] w_sys_tmp478;
	wire signed [31:0] w_sys_tmp659;
	wire               w_sys_tmp660;
	wire               w_sys_tmp661;
	wire signed [31:0] w_sys_tmp662;
	wire signed [31:0] w_sys_tmp665;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp667;
	wire        [31:0] w_sys_tmp668;
	wire signed [31:0] w_sys_tmp669;
	wire signed [31:0] w_sys_tmp670;
	wire signed [31:0] w_sys_tmp673;
	wire signed [31:0] w_sys_tmp674;
	wire        [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp677;
	wire signed [31:0] w_sys_tmp678;
	wire signed [31:0] w_sys_tmp681;
	wire signed [31:0] w_sys_tmp682;
	wire        [31:0] w_sys_tmp684;
	wire signed [31:0] w_sys_tmp685;
	wire signed [31:0] w_sys_tmp686;
	wire signed [31:0] w_sys_tmp688;
	wire signed [31:0] w_sys_tmp689;
	wire signed [31:0] w_sys_tmp690;
	wire signed [31:0] w_sys_tmp691;
	wire signed [31:0] w_sys_tmp692;
	wire signed [31:0] w_sys_tmp693;
	wire signed [31:0] w_sys_tmp874;
	wire               w_sys_tmp875;
	wire               w_sys_tmp876;
	wire signed [31:0] w_sys_tmp877;
	wire signed [31:0] w_sys_tmp880;
	wire signed [31:0] w_sys_tmp881;
	wire signed [31:0] w_sys_tmp882;
	wire        [31:0] w_sys_tmp883;
	wire signed [31:0] w_sys_tmp884;
	wire signed [31:0] w_sys_tmp885;
	wire signed [31:0] w_sys_tmp888;
	wire signed [31:0] w_sys_tmp889;
	wire        [31:0] w_sys_tmp891;
	wire signed [31:0] w_sys_tmp892;
	wire signed [31:0] w_sys_tmp893;
	wire signed [31:0] w_sys_tmp896;
	wire signed [31:0] w_sys_tmp897;
	wire        [31:0] w_sys_tmp899;
	wire signed [31:0] w_sys_tmp900;
	wire signed [31:0] w_sys_tmp901;
	wire signed [31:0] w_sys_tmp903;
	wire signed [31:0] w_sys_tmp904;
	wire signed [31:0] w_sys_tmp905;
	wire signed [31:0] w_sys_tmp906;
	wire signed [31:0] w_sys_tmp907;
	wire signed [31:0] w_sys_tmp908;
	wire signed [31:0] w_sys_tmp1089;
	wire               w_sys_tmp1090;
	wire               w_sys_tmp1091;
	wire signed [31:0] w_sys_tmp1092;
	wire signed [31:0] w_sys_tmp1095;
	wire signed [31:0] w_sys_tmp1096;
	wire signed [31:0] w_sys_tmp1097;
	wire        [31:0] w_sys_tmp1098;
	wire signed [31:0] w_sys_tmp1099;
	wire signed [31:0] w_sys_tmp1100;
	wire signed [31:0] w_sys_tmp1103;
	wire signed [31:0] w_sys_tmp1104;
	wire        [31:0] w_sys_tmp1106;
	wire signed [31:0] w_sys_tmp1107;
	wire signed [31:0] w_sys_tmp1108;
	wire signed [31:0] w_sys_tmp1111;
	wire signed [31:0] w_sys_tmp1112;
	wire        [31:0] w_sys_tmp1114;
	wire signed [31:0] w_sys_tmp1115;
	wire signed [31:0] w_sys_tmp1116;
	wire signed [31:0] w_sys_tmp1118;
	wire signed [31:0] w_sys_tmp1119;
	wire signed [31:0] w_sys_tmp1120;
	wire signed [31:0] w_sys_tmp1121;
	wire signed [31:0] w_sys_tmp1122;
	wire signed [31:0] w_sys_tmp1123;
	wire signed [31:0] w_sys_tmp1304;
	wire               w_sys_tmp1305;
	wire               w_sys_tmp1306;
	wire signed [31:0] w_sys_tmp1307;
	wire signed [31:0] w_sys_tmp1310;
	wire signed [31:0] w_sys_tmp1311;
	wire signed [31:0] w_sys_tmp1312;
	wire        [31:0] w_sys_tmp1313;
	wire signed [31:0] w_sys_tmp1314;
	wire signed [31:0] w_sys_tmp1315;
	wire signed [31:0] w_sys_tmp1318;
	wire signed [31:0] w_sys_tmp1319;
	wire        [31:0] w_sys_tmp1321;
	wire signed [31:0] w_sys_tmp1322;
	wire signed [31:0] w_sys_tmp1323;
	wire signed [31:0] w_sys_tmp1326;
	wire signed [31:0] w_sys_tmp1327;
	wire        [31:0] w_sys_tmp1329;
	wire signed [31:0] w_sys_tmp1330;
	wire signed [31:0] w_sys_tmp1331;
	wire signed [31:0] w_sys_tmp1333;
	wire signed [31:0] w_sys_tmp1334;
	wire signed [31:0] w_sys_tmp1335;
	wire signed [31:0] w_sys_tmp1336;
	wire signed [31:0] w_sys_tmp1337;
	wire signed [31:0] w_sys_tmp1338;
	wire signed [31:0] w_sys_tmp1519;
	wire               w_sys_tmp1520;
	wire               w_sys_tmp1521;
	wire signed [31:0] w_sys_tmp1522;
	wire signed [31:0] w_sys_tmp1525;
	wire signed [31:0] w_sys_tmp1526;
	wire signed [31:0] w_sys_tmp1527;
	wire        [31:0] w_sys_tmp1528;
	wire signed [31:0] w_sys_tmp1529;
	wire signed [31:0] w_sys_tmp1530;
	wire signed [31:0] w_sys_tmp1533;
	wire signed [31:0] w_sys_tmp1534;
	wire        [31:0] w_sys_tmp1536;
	wire signed [31:0] w_sys_tmp1537;
	wire signed [31:0] w_sys_tmp1538;
	wire signed [31:0] w_sys_tmp1541;
	wire signed [31:0] w_sys_tmp1542;
	wire        [31:0] w_sys_tmp1544;
	wire signed [31:0] w_sys_tmp1545;
	wire signed [31:0] w_sys_tmp1546;
	wire signed [31:0] w_sys_tmp1548;
	wire signed [31:0] w_sys_tmp1549;
	wire signed [31:0] w_sys_tmp1550;
	wire signed [31:0] w_sys_tmp1551;
	wire signed [31:0] w_sys_tmp1552;
	wire signed [31:0] w_sys_tmp1553;
	wire signed [31:0] w_sys_tmp1734;
	wire               w_sys_tmp1735;
	wire               w_sys_tmp1736;
	wire signed [31:0] w_sys_tmp1737;
	wire signed [31:0] w_sys_tmp1740;
	wire signed [31:0] w_sys_tmp1741;
	wire signed [31:0] w_sys_tmp1742;
	wire        [31:0] w_sys_tmp1743;
	wire signed [31:0] w_sys_tmp1744;
	wire signed [31:0] w_sys_tmp1745;
	wire signed [31:0] w_sys_tmp1748;
	wire signed [31:0] w_sys_tmp1749;
	wire        [31:0] w_sys_tmp1751;
	wire signed [31:0] w_sys_tmp1752;
	wire signed [31:0] w_sys_tmp1753;
	wire signed [31:0] w_sys_tmp1756;
	wire signed [31:0] w_sys_tmp1757;
	wire        [31:0] w_sys_tmp1759;
	wire signed [31:0] w_sys_tmp1760;
	wire signed [31:0] w_sys_tmp1761;
	wire signed [31:0] w_sys_tmp1763;
	wire signed [31:0] w_sys_tmp1764;
	wire signed [31:0] w_sys_tmp1765;
	wire signed [31:0] w_sys_tmp1766;
	wire signed [31:0] w_sys_tmp1767;
	wire signed [31:0] w_sys_tmp1768;
	wire               w_sys_tmp1949;
	wire               w_sys_tmp1950;
	wire signed [31:0] w_sys_tmp1951;
	wire signed [31:0] w_sys_tmp1952;
	wire               w_sys_tmp1953;
	wire               w_sys_tmp1954;
	wire signed [31:0] w_sys_tmp1955;
	wire signed [31:0] w_sys_tmp1958;
	wire signed [31:0] w_sys_tmp1959;
	wire signed [31:0] w_sys_tmp1960;
	wire        [31:0] w_sys_tmp1961;
	wire signed [31:0] w_sys_tmp1962;
	wire signed [31:0] w_sys_tmp1963;
	wire signed [31:0] w_sys_tmp1966;
	wire signed [31:0] w_sys_tmp1967;
	wire        [31:0] w_sys_tmp1969;
	wire signed [31:0] w_sys_tmp1970;
	wire signed [31:0] w_sys_tmp1971;
	wire signed [31:0] w_sys_tmp1974;
	wire signed [31:0] w_sys_tmp1975;
	wire        [31:0] w_sys_tmp1977;
	wire signed [31:0] w_sys_tmp1978;
	wire signed [31:0] w_sys_tmp1979;
	wire signed [31:0] w_sys_tmp1981;
	wire signed [31:0] w_sys_tmp1982;
	wire signed [31:0] w_sys_tmp1983;
	wire signed [31:0] w_sys_tmp1984;
	wire signed [31:0] w_sys_tmp1985;
	wire signed [31:0] w_sys_tmp1986;
	wire signed [31:0] w_sys_tmp2167;
	wire               w_sys_tmp2168;
	wire               w_sys_tmp2169;
	wire signed [31:0] w_sys_tmp2170;
	wire signed [31:0] w_sys_tmp2173;
	wire signed [31:0] w_sys_tmp2174;
	wire signed [31:0] w_sys_tmp2175;
	wire        [31:0] w_sys_tmp2176;
	wire signed [31:0] w_sys_tmp2177;
	wire signed [31:0] w_sys_tmp2178;
	wire signed [31:0] w_sys_tmp2181;
	wire signed [31:0] w_sys_tmp2182;
	wire        [31:0] w_sys_tmp2184;
	wire signed [31:0] w_sys_tmp2185;
	wire signed [31:0] w_sys_tmp2186;
	wire signed [31:0] w_sys_tmp2189;
	wire signed [31:0] w_sys_tmp2190;
	wire        [31:0] w_sys_tmp2192;
	wire signed [31:0] w_sys_tmp2193;
	wire signed [31:0] w_sys_tmp2194;
	wire signed [31:0] w_sys_tmp2196;
	wire signed [31:0] w_sys_tmp2197;
	wire signed [31:0] w_sys_tmp2198;
	wire signed [31:0] w_sys_tmp2199;
	wire signed [31:0] w_sys_tmp2200;
	wire signed [31:0] w_sys_tmp2201;
	wire signed [31:0] w_sys_tmp2382;
	wire               w_sys_tmp2383;
	wire               w_sys_tmp2384;
	wire signed [31:0] w_sys_tmp2385;
	wire signed [31:0] w_sys_tmp2388;
	wire signed [31:0] w_sys_tmp2389;
	wire signed [31:0] w_sys_tmp2390;
	wire        [31:0] w_sys_tmp2391;
	wire signed [31:0] w_sys_tmp2392;
	wire signed [31:0] w_sys_tmp2393;
	wire signed [31:0] w_sys_tmp2396;
	wire signed [31:0] w_sys_tmp2397;
	wire        [31:0] w_sys_tmp2399;
	wire signed [31:0] w_sys_tmp2400;
	wire signed [31:0] w_sys_tmp2401;
	wire signed [31:0] w_sys_tmp2404;
	wire signed [31:0] w_sys_tmp2405;
	wire        [31:0] w_sys_tmp2407;
	wire signed [31:0] w_sys_tmp2408;
	wire signed [31:0] w_sys_tmp2409;
	wire signed [31:0] w_sys_tmp2411;
	wire signed [31:0] w_sys_tmp2412;
	wire signed [31:0] w_sys_tmp2413;
	wire signed [31:0] w_sys_tmp2414;
	wire signed [31:0] w_sys_tmp2415;
	wire signed [31:0] w_sys_tmp2416;
	wire signed [31:0] w_sys_tmp2597;
	wire               w_sys_tmp2598;
	wire               w_sys_tmp2599;
	wire signed [31:0] w_sys_tmp2600;
	wire signed [31:0] w_sys_tmp2603;
	wire signed [31:0] w_sys_tmp2604;
	wire signed [31:0] w_sys_tmp2605;
	wire        [31:0] w_sys_tmp2606;
	wire signed [31:0] w_sys_tmp2607;
	wire signed [31:0] w_sys_tmp2608;
	wire signed [31:0] w_sys_tmp2611;
	wire signed [31:0] w_sys_tmp2612;
	wire        [31:0] w_sys_tmp2614;
	wire signed [31:0] w_sys_tmp2615;
	wire signed [31:0] w_sys_tmp2616;
	wire signed [31:0] w_sys_tmp2619;
	wire signed [31:0] w_sys_tmp2620;
	wire        [31:0] w_sys_tmp2622;
	wire signed [31:0] w_sys_tmp2623;
	wire signed [31:0] w_sys_tmp2624;
	wire signed [31:0] w_sys_tmp2626;
	wire signed [31:0] w_sys_tmp2627;
	wire signed [31:0] w_sys_tmp2628;
	wire signed [31:0] w_sys_tmp2629;
	wire signed [31:0] w_sys_tmp2630;
	wire signed [31:0] w_sys_tmp2631;
	wire signed [31:0] w_sys_tmp2812;
	wire               w_sys_tmp2813;
	wire               w_sys_tmp2814;
	wire signed [31:0] w_sys_tmp2815;
	wire signed [31:0] w_sys_tmp2818;
	wire signed [31:0] w_sys_tmp2819;
	wire signed [31:0] w_sys_tmp2820;
	wire        [31:0] w_sys_tmp2821;
	wire signed [31:0] w_sys_tmp2822;
	wire signed [31:0] w_sys_tmp2823;
	wire signed [31:0] w_sys_tmp2826;
	wire signed [31:0] w_sys_tmp2827;
	wire        [31:0] w_sys_tmp2829;
	wire signed [31:0] w_sys_tmp2830;
	wire signed [31:0] w_sys_tmp2831;
	wire signed [31:0] w_sys_tmp2834;
	wire signed [31:0] w_sys_tmp2835;
	wire        [31:0] w_sys_tmp2837;
	wire signed [31:0] w_sys_tmp2838;
	wire signed [31:0] w_sys_tmp2839;
	wire signed [31:0] w_sys_tmp2841;
	wire signed [31:0] w_sys_tmp2842;
	wire signed [31:0] w_sys_tmp2843;
	wire signed [31:0] w_sys_tmp2844;
	wire signed [31:0] w_sys_tmp2845;
	wire signed [31:0] w_sys_tmp2846;
	wire signed [31:0] w_sys_tmp3027;
	wire               w_sys_tmp3028;
	wire               w_sys_tmp3029;
	wire signed [31:0] w_sys_tmp3030;
	wire signed [31:0] w_sys_tmp3033;
	wire signed [31:0] w_sys_tmp3034;
	wire signed [31:0] w_sys_tmp3035;
	wire        [31:0] w_sys_tmp3036;
	wire signed [31:0] w_sys_tmp3037;
	wire signed [31:0] w_sys_tmp3038;
	wire signed [31:0] w_sys_tmp3041;
	wire signed [31:0] w_sys_tmp3042;
	wire        [31:0] w_sys_tmp3044;
	wire signed [31:0] w_sys_tmp3045;
	wire signed [31:0] w_sys_tmp3046;
	wire signed [31:0] w_sys_tmp3049;
	wire signed [31:0] w_sys_tmp3050;
	wire        [31:0] w_sys_tmp3052;
	wire signed [31:0] w_sys_tmp3053;
	wire signed [31:0] w_sys_tmp3054;
	wire signed [31:0] w_sys_tmp3056;
	wire signed [31:0] w_sys_tmp3057;
	wire signed [31:0] w_sys_tmp3058;
	wire signed [31:0] w_sys_tmp3059;
	wire signed [31:0] w_sys_tmp3060;
	wire signed [31:0] w_sys_tmp3061;
	wire signed [31:0] w_sys_tmp3242;
	wire               w_sys_tmp3243;
	wire               w_sys_tmp3244;
	wire signed [31:0] w_sys_tmp3245;
	wire signed [31:0] w_sys_tmp3248;
	wire signed [31:0] w_sys_tmp3249;
	wire signed [31:0] w_sys_tmp3250;
	wire        [31:0] w_sys_tmp3251;
	wire signed [31:0] w_sys_tmp3252;
	wire signed [31:0] w_sys_tmp3253;
	wire signed [31:0] w_sys_tmp3256;
	wire signed [31:0] w_sys_tmp3257;
	wire        [31:0] w_sys_tmp3259;
	wire signed [31:0] w_sys_tmp3260;
	wire signed [31:0] w_sys_tmp3261;
	wire signed [31:0] w_sys_tmp3264;
	wire signed [31:0] w_sys_tmp3265;
	wire        [31:0] w_sys_tmp3267;
	wire signed [31:0] w_sys_tmp3268;
	wire signed [31:0] w_sys_tmp3269;
	wire signed [31:0] w_sys_tmp3271;
	wire signed [31:0] w_sys_tmp3272;
	wire signed [31:0] w_sys_tmp3273;
	wire signed [31:0] w_sys_tmp3274;
	wire signed [31:0] w_sys_tmp3275;
	wire signed [31:0] w_sys_tmp3276;
	wire signed [31:0] w_sys_tmp3457;
	wire               w_sys_tmp3458;
	wire               w_sys_tmp3459;
	wire signed [31:0] w_sys_tmp3460;
	wire signed [31:0] w_sys_tmp3463;
	wire signed [31:0] w_sys_tmp3464;
	wire signed [31:0] w_sys_tmp3465;
	wire        [31:0] w_sys_tmp3466;
	wire signed [31:0] w_sys_tmp3467;
	wire signed [31:0] w_sys_tmp3468;
	wire signed [31:0] w_sys_tmp3471;
	wire signed [31:0] w_sys_tmp3472;
	wire        [31:0] w_sys_tmp3474;
	wire signed [31:0] w_sys_tmp3475;
	wire signed [31:0] w_sys_tmp3476;
	wire signed [31:0] w_sys_tmp3479;
	wire signed [31:0] w_sys_tmp3480;
	wire        [31:0] w_sys_tmp3482;
	wire signed [31:0] w_sys_tmp3483;
	wire signed [31:0] w_sys_tmp3484;
	wire signed [31:0] w_sys_tmp3486;
	wire signed [31:0] w_sys_tmp3487;
	wire signed [31:0] w_sys_tmp3488;
	wire signed [31:0] w_sys_tmp3489;
	wire signed [31:0] w_sys_tmp3490;
	wire signed [31:0] w_sys_tmp3491;
	wire               w_sys_tmp3672;
	wire               w_sys_tmp3673;
	wire signed [31:0] w_sys_tmp3674;
	wire signed [31:0] w_sys_tmp3675;
	wire               w_sys_tmp3676;
	wire               w_sys_tmp3677;
	wire signed [31:0] w_sys_tmp3678;
	wire signed [31:0] w_sys_tmp3681;
	wire signed [31:0] w_sys_tmp3682;
	wire signed [31:0] w_sys_tmp3683;
	wire        [31:0] w_sys_tmp3684;
	wire signed [31:0] w_sys_tmp3685;
	wire signed [31:0] w_sys_tmp3686;
	wire signed [31:0] w_sys_tmp3689;
	wire signed [31:0] w_sys_tmp3690;
	wire        [31:0] w_sys_tmp3692;
	wire signed [31:0] w_sys_tmp3693;
	wire signed [31:0] w_sys_tmp3694;
	wire signed [31:0] w_sys_tmp3697;
	wire signed [31:0] w_sys_tmp3698;
	wire        [31:0] w_sys_tmp3700;
	wire signed [31:0] w_sys_tmp3701;
	wire signed [31:0] w_sys_tmp3702;
	wire signed [31:0] w_sys_tmp3704;
	wire signed [31:0] w_sys_tmp3705;
	wire signed [31:0] w_sys_tmp3706;
	wire signed [31:0] w_sys_tmp3707;
	wire signed [31:0] w_sys_tmp3708;
	wire signed [31:0] w_sys_tmp3709;
	wire signed [31:0] w_sys_tmp3890;
	wire               w_sys_tmp3891;
	wire               w_sys_tmp3892;
	wire signed [31:0] w_sys_tmp3893;
	wire signed [31:0] w_sys_tmp3896;
	wire signed [31:0] w_sys_tmp3897;
	wire signed [31:0] w_sys_tmp3898;
	wire        [31:0] w_sys_tmp3899;
	wire signed [31:0] w_sys_tmp3900;
	wire signed [31:0] w_sys_tmp3901;
	wire signed [31:0] w_sys_tmp3904;
	wire signed [31:0] w_sys_tmp3905;
	wire        [31:0] w_sys_tmp3907;
	wire signed [31:0] w_sys_tmp3908;
	wire signed [31:0] w_sys_tmp3909;
	wire signed [31:0] w_sys_tmp3912;
	wire signed [31:0] w_sys_tmp3913;
	wire        [31:0] w_sys_tmp3915;
	wire signed [31:0] w_sys_tmp3916;
	wire signed [31:0] w_sys_tmp3917;
	wire signed [31:0] w_sys_tmp3919;
	wire signed [31:0] w_sys_tmp3920;
	wire signed [31:0] w_sys_tmp3921;
	wire signed [31:0] w_sys_tmp3922;
	wire signed [31:0] w_sys_tmp3923;
	wire signed [31:0] w_sys_tmp3924;
	wire signed [31:0] w_sys_tmp4105;
	wire               w_sys_tmp4106;
	wire               w_sys_tmp4107;
	wire signed [31:0] w_sys_tmp4108;
	wire signed [31:0] w_sys_tmp4111;
	wire signed [31:0] w_sys_tmp4112;
	wire signed [31:0] w_sys_tmp4113;
	wire        [31:0] w_sys_tmp4114;
	wire signed [31:0] w_sys_tmp4115;
	wire signed [31:0] w_sys_tmp4116;
	wire signed [31:0] w_sys_tmp4119;
	wire signed [31:0] w_sys_tmp4120;
	wire        [31:0] w_sys_tmp4122;
	wire signed [31:0] w_sys_tmp4123;
	wire signed [31:0] w_sys_tmp4124;
	wire signed [31:0] w_sys_tmp4127;
	wire signed [31:0] w_sys_tmp4128;
	wire        [31:0] w_sys_tmp4130;
	wire signed [31:0] w_sys_tmp4131;
	wire signed [31:0] w_sys_tmp4132;
	wire signed [31:0] w_sys_tmp4134;
	wire signed [31:0] w_sys_tmp4135;
	wire signed [31:0] w_sys_tmp4136;
	wire signed [31:0] w_sys_tmp4137;
	wire signed [31:0] w_sys_tmp4138;
	wire signed [31:0] w_sys_tmp4139;
	wire signed [31:0] w_sys_tmp4320;
	wire               w_sys_tmp4321;
	wire               w_sys_tmp4322;
	wire signed [31:0] w_sys_tmp4323;
	wire signed [31:0] w_sys_tmp4326;
	wire signed [31:0] w_sys_tmp4327;
	wire signed [31:0] w_sys_tmp4328;
	wire        [31:0] w_sys_tmp4329;
	wire signed [31:0] w_sys_tmp4330;
	wire signed [31:0] w_sys_tmp4331;
	wire signed [31:0] w_sys_tmp4334;
	wire signed [31:0] w_sys_tmp4335;
	wire        [31:0] w_sys_tmp4337;
	wire signed [31:0] w_sys_tmp4338;
	wire signed [31:0] w_sys_tmp4339;
	wire signed [31:0] w_sys_tmp4342;
	wire signed [31:0] w_sys_tmp4343;
	wire        [31:0] w_sys_tmp4345;
	wire signed [31:0] w_sys_tmp4346;
	wire signed [31:0] w_sys_tmp4347;
	wire signed [31:0] w_sys_tmp4349;
	wire signed [31:0] w_sys_tmp4350;
	wire signed [31:0] w_sys_tmp4351;
	wire signed [31:0] w_sys_tmp4352;
	wire signed [31:0] w_sys_tmp4353;
	wire signed [31:0] w_sys_tmp4354;
	wire signed [31:0] w_sys_tmp4535;
	wire               w_sys_tmp4536;
	wire               w_sys_tmp4537;
	wire signed [31:0] w_sys_tmp4538;
	wire signed [31:0] w_sys_tmp4541;
	wire signed [31:0] w_sys_tmp4542;
	wire signed [31:0] w_sys_tmp4543;
	wire        [31:0] w_sys_tmp4544;
	wire signed [31:0] w_sys_tmp4545;
	wire signed [31:0] w_sys_tmp4546;
	wire signed [31:0] w_sys_tmp4549;
	wire signed [31:0] w_sys_tmp4550;
	wire        [31:0] w_sys_tmp4552;
	wire signed [31:0] w_sys_tmp4553;
	wire signed [31:0] w_sys_tmp4554;
	wire signed [31:0] w_sys_tmp4557;
	wire signed [31:0] w_sys_tmp4558;
	wire        [31:0] w_sys_tmp4560;
	wire signed [31:0] w_sys_tmp4561;
	wire signed [31:0] w_sys_tmp4562;
	wire signed [31:0] w_sys_tmp4564;
	wire signed [31:0] w_sys_tmp4565;
	wire signed [31:0] w_sys_tmp4566;
	wire signed [31:0] w_sys_tmp4567;
	wire signed [31:0] w_sys_tmp4568;
	wire signed [31:0] w_sys_tmp4569;
	wire signed [31:0] w_sys_tmp4750;
	wire               w_sys_tmp4751;
	wire               w_sys_tmp4752;
	wire signed [31:0] w_sys_tmp4753;
	wire signed [31:0] w_sys_tmp4756;
	wire signed [31:0] w_sys_tmp4757;
	wire signed [31:0] w_sys_tmp4758;
	wire        [31:0] w_sys_tmp4759;
	wire signed [31:0] w_sys_tmp4760;
	wire signed [31:0] w_sys_tmp4761;
	wire signed [31:0] w_sys_tmp4764;
	wire signed [31:0] w_sys_tmp4765;
	wire        [31:0] w_sys_tmp4767;
	wire signed [31:0] w_sys_tmp4768;
	wire signed [31:0] w_sys_tmp4769;
	wire signed [31:0] w_sys_tmp4772;
	wire signed [31:0] w_sys_tmp4773;
	wire        [31:0] w_sys_tmp4775;
	wire signed [31:0] w_sys_tmp4776;
	wire signed [31:0] w_sys_tmp4777;
	wire signed [31:0] w_sys_tmp4779;
	wire signed [31:0] w_sys_tmp4780;
	wire signed [31:0] w_sys_tmp4781;
	wire signed [31:0] w_sys_tmp4782;
	wire signed [31:0] w_sys_tmp4783;
	wire signed [31:0] w_sys_tmp4784;
	wire signed [31:0] w_sys_tmp4965;
	wire               w_sys_tmp4966;
	wire               w_sys_tmp4967;
	wire signed [31:0] w_sys_tmp4968;
	wire signed [31:0] w_sys_tmp4971;
	wire signed [31:0] w_sys_tmp4972;
	wire signed [31:0] w_sys_tmp4973;
	wire        [31:0] w_sys_tmp4974;
	wire signed [31:0] w_sys_tmp4975;
	wire signed [31:0] w_sys_tmp4976;
	wire signed [31:0] w_sys_tmp4979;
	wire signed [31:0] w_sys_tmp4980;
	wire        [31:0] w_sys_tmp4982;
	wire signed [31:0] w_sys_tmp4983;
	wire signed [31:0] w_sys_tmp4984;
	wire signed [31:0] w_sys_tmp4987;
	wire signed [31:0] w_sys_tmp4988;
	wire        [31:0] w_sys_tmp4990;
	wire signed [31:0] w_sys_tmp4991;
	wire signed [31:0] w_sys_tmp4992;
	wire signed [31:0] w_sys_tmp4994;
	wire signed [31:0] w_sys_tmp4995;
	wire signed [31:0] w_sys_tmp4996;
	wire signed [31:0] w_sys_tmp4997;
	wire signed [31:0] w_sys_tmp4998;
	wire signed [31:0] w_sys_tmp4999;
	wire signed [31:0] w_sys_tmp5180;
	wire               w_sys_tmp5181;
	wire               w_sys_tmp5182;
	wire signed [31:0] w_sys_tmp5183;
	wire signed [31:0] w_sys_tmp5186;
	wire signed [31:0] w_sys_tmp5187;
	wire signed [31:0] w_sys_tmp5188;
	wire        [31:0] w_sys_tmp5189;
	wire signed [31:0] w_sys_tmp5190;
	wire signed [31:0] w_sys_tmp5191;
	wire signed [31:0] w_sys_tmp5194;
	wire signed [31:0] w_sys_tmp5195;
	wire        [31:0] w_sys_tmp5197;
	wire signed [31:0] w_sys_tmp5198;
	wire signed [31:0] w_sys_tmp5199;
	wire signed [31:0] w_sys_tmp5202;
	wire signed [31:0] w_sys_tmp5203;
	wire        [31:0] w_sys_tmp5205;
	wire signed [31:0] w_sys_tmp5206;
	wire signed [31:0] w_sys_tmp5207;
	wire signed [31:0] w_sys_tmp5209;
	wire signed [31:0] w_sys_tmp5210;
	wire signed [31:0] w_sys_tmp5211;
	wire signed [31:0] w_sys_tmp5212;
	wire signed [31:0] w_sys_tmp5213;
	wire signed [31:0] w_sys_tmp5214;
	wire               w_sys_tmp5395;
	wire               w_sys_tmp5396;
	wire signed [31:0] w_sys_tmp5397;
	wire signed [31:0] w_sys_tmp5398;
	wire               w_sys_tmp5399;
	wire               w_sys_tmp5400;
	wire signed [31:0] w_sys_tmp5401;
	wire signed [31:0] w_sys_tmp5404;
	wire signed [31:0] w_sys_tmp5405;
	wire signed [31:0] w_sys_tmp5406;
	wire        [31:0] w_sys_tmp5407;
	wire signed [31:0] w_sys_tmp5408;
	wire signed [31:0] w_sys_tmp5409;
	wire signed [31:0] w_sys_tmp5412;
	wire signed [31:0] w_sys_tmp5413;
	wire        [31:0] w_sys_tmp5415;
	wire signed [31:0] w_sys_tmp5416;
	wire signed [31:0] w_sys_tmp5417;
	wire signed [31:0] w_sys_tmp5420;
	wire signed [31:0] w_sys_tmp5421;
	wire        [31:0] w_sys_tmp5423;
	wire signed [31:0] w_sys_tmp5424;
	wire signed [31:0] w_sys_tmp5425;
	wire signed [31:0] w_sys_tmp5427;
	wire signed [31:0] w_sys_tmp5428;
	wire signed [31:0] w_sys_tmp5429;
	wire signed [31:0] w_sys_tmp5430;
	wire signed [31:0] w_sys_tmp5431;
	wire signed [31:0] w_sys_tmp5432;
	wire signed [31:0] w_sys_tmp5613;
	wire               w_sys_tmp5614;
	wire               w_sys_tmp5615;
	wire signed [31:0] w_sys_tmp5616;
	wire signed [31:0] w_sys_tmp5619;
	wire signed [31:0] w_sys_tmp5620;
	wire signed [31:0] w_sys_tmp5621;
	wire        [31:0] w_sys_tmp5622;
	wire signed [31:0] w_sys_tmp5623;
	wire signed [31:0] w_sys_tmp5624;
	wire signed [31:0] w_sys_tmp5627;
	wire signed [31:0] w_sys_tmp5628;
	wire        [31:0] w_sys_tmp5630;
	wire signed [31:0] w_sys_tmp5631;
	wire signed [31:0] w_sys_tmp5632;
	wire signed [31:0] w_sys_tmp5635;
	wire signed [31:0] w_sys_tmp5636;
	wire        [31:0] w_sys_tmp5638;
	wire signed [31:0] w_sys_tmp5639;
	wire signed [31:0] w_sys_tmp5640;
	wire signed [31:0] w_sys_tmp5642;
	wire signed [31:0] w_sys_tmp5643;
	wire signed [31:0] w_sys_tmp5644;
	wire signed [31:0] w_sys_tmp5645;
	wire signed [31:0] w_sys_tmp5646;
	wire signed [31:0] w_sys_tmp5647;
	wire signed [31:0] w_sys_tmp5828;
	wire               w_sys_tmp5829;
	wire               w_sys_tmp5830;
	wire signed [31:0] w_sys_tmp5831;
	wire signed [31:0] w_sys_tmp5834;
	wire signed [31:0] w_sys_tmp5835;
	wire signed [31:0] w_sys_tmp5836;
	wire        [31:0] w_sys_tmp5837;
	wire signed [31:0] w_sys_tmp5838;
	wire signed [31:0] w_sys_tmp5839;
	wire signed [31:0] w_sys_tmp5842;
	wire signed [31:0] w_sys_tmp5843;
	wire        [31:0] w_sys_tmp5845;
	wire signed [31:0] w_sys_tmp5846;
	wire signed [31:0] w_sys_tmp5847;
	wire signed [31:0] w_sys_tmp5850;
	wire signed [31:0] w_sys_tmp5851;
	wire        [31:0] w_sys_tmp5853;
	wire signed [31:0] w_sys_tmp5854;
	wire signed [31:0] w_sys_tmp5855;
	wire signed [31:0] w_sys_tmp5857;
	wire signed [31:0] w_sys_tmp5858;
	wire signed [31:0] w_sys_tmp5859;
	wire signed [31:0] w_sys_tmp5860;
	wire signed [31:0] w_sys_tmp5861;
	wire signed [31:0] w_sys_tmp5862;
	wire signed [31:0] w_sys_tmp6043;
	wire               w_sys_tmp6044;
	wire               w_sys_tmp6045;
	wire signed [31:0] w_sys_tmp6046;
	wire signed [31:0] w_sys_tmp6049;
	wire signed [31:0] w_sys_tmp6050;
	wire signed [31:0] w_sys_tmp6051;
	wire        [31:0] w_sys_tmp6052;
	wire signed [31:0] w_sys_tmp6053;
	wire signed [31:0] w_sys_tmp6054;
	wire signed [31:0] w_sys_tmp6057;
	wire signed [31:0] w_sys_tmp6058;
	wire        [31:0] w_sys_tmp6060;
	wire signed [31:0] w_sys_tmp6061;
	wire signed [31:0] w_sys_tmp6062;
	wire signed [31:0] w_sys_tmp6065;
	wire signed [31:0] w_sys_tmp6066;
	wire        [31:0] w_sys_tmp6068;
	wire signed [31:0] w_sys_tmp6069;
	wire signed [31:0] w_sys_tmp6070;
	wire signed [31:0] w_sys_tmp6072;
	wire signed [31:0] w_sys_tmp6073;
	wire signed [31:0] w_sys_tmp6074;
	wire signed [31:0] w_sys_tmp6075;
	wire signed [31:0] w_sys_tmp6076;
	wire signed [31:0] w_sys_tmp6077;
	wire signed [31:0] w_sys_tmp6258;
	wire               w_sys_tmp6259;
	wire               w_sys_tmp6260;
	wire signed [31:0] w_sys_tmp6261;
	wire signed [31:0] w_sys_tmp6264;
	wire signed [31:0] w_sys_tmp6265;
	wire signed [31:0] w_sys_tmp6266;
	wire        [31:0] w_sys_tmp6267;
	wire signed [31:0] w_sys_tmp6268;
	wire signed [31:0] w_sys_tmp6269;
	wire signed [31:0] w_sys_tmp6272;
	wire signed [31:0] w_sys_tmp6273;
	wire        [31:0] w_sys_tmp6275;
	wire signed [31:0] w_sys_tmp6276;
	wire signed [31:0] w_sys_tmp6277;
	wire signed [31:0] w_sys_tmp6280;
	wire signed [31:0] w_sys_tmp6281;
	wire        [31:0] w_sys_tmp6283;
	wire signed [31:0] w_sys_tmp6284;
	wire signed [31:0] w_sys_tmp6285;
	wire signed [31:0] w_sys_tmp6287;
	wire signed [31:0] w_sys_tmp6288;
	wire signed [31:0] w_sys_tmp6289;
	wire signed [31:0] w_sys_tmp6290;
	wire signed [31:0] w_sys_tmp6291;
	wire signed [31:0] w_sys_tmp6292;
	wire signed [31:0] w_sys_tmp6473;
	wire               w_sys_tmp6474;
	wire               w_sys_tmp6475;
	wire signed [31:0] w_sys_tmp6476;
	wire signed [31:0] w_sys_tmp6479;
	wire signed [31:0] w_sys_tmp6480;
	wire signed [31:0] w_sys_tmp6481;
	wire        [31:0] w_sys_tmp6482;
	wire signed [31:0] w_sys_tmp6483;
	wire signed [31:0] w_sys_tmp6484;
	wire signed [31:0] w_sys_tmp6487;
	wire signed [31:0] w_sys_tmp6488;
	wire        [31:0] w_sys_tmp6490;
	wire signed [31:0] w_sys_tmp6491;
	wire signed [31:0] w_sys_tmp6492;
	wire signed [31:0] w_sys_tmp6495;
	wire signed [31:0] w_sys_tmp6496;
	wire        [31:0] w_sys_tmp6498;
	wire signed [31:0] w_sys_tmp6499;
	wire signed [31:0] w_sys_tmp6500;
	wire signed [31:0] w_sys_tmp6502;
	wire signed [31:0] w_sys_tmp6503;
	wire signed [31:0] w_sys_tmp6504;
	wire signed [31:0] w_sys_tmp6505;
	wire signed [31:0] w_sys_tmp6506;
	wire signed [31:0] w_sys_tmp6507;
	wire signed [31:0] w_sys_tmp6688;
	wire               w_sys_tmp6689;
	wire               w_sys_tmp6690;
	wire signed [31:0] w_sys_tmp6691;
	wire signed [31:0] w_sys_tmp6694;
	wire signed [31:0] w_sys_tmp6695;
	wire signed [31:0] w_sys_tmp6696;
	wire        [31:0] w_sys_tmp6697;
	wire signed [31:0] w_sys_tmp6698;
	wire signed [31:0] w_sys_tmp6699;
	wire signed [31:0] w_sys_tmp6702;
	wire signed [31:0] w_sys_tmp6703;
	wire        [31:0] w_sys_tmp6705;
	wire signed [31:0] w_sys_tmp6706;
	wire signed [31:0] w_sys_tmp6707;
	wire signed [31:0] w_sys_tmp6710;
	wire signed [31:0] w_sys_tmp6711;
	wire        [31:0] w_sys_tmp6713;
	wire signed [31:0] w_sys_tmp6714;
	wire signed [31:0] w_sys_tmp6715;
	wire signed [31:0] w_sys_tmp6717;
	wire signed [31:0] w_sys_tmp6718;
	wire signed [31:0] w_sys_tmp6719;
	wire signed [31:0] w_sys_tmp6720;
	wire signed [31:0] w_sys_tmp6721;
	wire signed [31:0] w_sys_tmp6722;
	wire signed [31:0] w_sys_tmp6903;
	wire               w_sys_tmp6904;
	wire               w_sys_tmp6905;
	wire signed [31:0] w_sys_tmp6906;
	wire signed [31:0] w_sys_tmp6909;
	wire signed [31:0] w_sys_tmp6910;
	wire signed [31:0] w_sys_tmp6911;
	wire        [31:0] w_sys_tmp6912;
	wire signed [31:0] w_sys_tmp6913;
	wire signed [31:0] w_sys_tmp6914;
	wire signed [31:0] w_sys_tmp6917;
	wire signed [31:0] w_sys_tmp6918;
	wire        [31:0] w_sys_tmp6920;
	wire signed [31:0] w_sys_tmp6921;
	wire signed [31:0] w_sys_tmp6922;
	wire signed [31:0] w_sys_tmp6925;
	wire signed [31:0] w_sys_tmp6926;
	wire        [31:0] w_sys_tmp6928;
	wire signed [31:0] w_sys_tmp6929;
	wire signed [31:0] w_sys_tmp6930;
	wire signed [31:0] w_sys_tmp6932;
	wire signed [31:0] w_sys_tmp6933;
	wire signed [31:0] w_sys_tmp6934;
	wire signed [31:0] w_sys_tmp6935;
	wire signed [31:0] w_sys_tmp6936;
	wire signed [31:0] w_sys_tmp6937;
	wire               w_sys_tmp7118;
	wire               w_sys_tmp7119;
	wire signed [31:0] w_sys_tmp7120;
	wire signed [31:0] w_sys_tmp7121;
	wire               w_sys_tmp7122;
	wire               w_sys_tmp7123;
	wire signed [31:0] w_sys_tmp7124;
	wire signed [31:0] w_sys_tmp7127;
	wire signed [31:0] w_sys_tmp7128;
	wire        [31:0] w_sys_tmp7129;
	wire signed [31:0] w_sys_tmp7130;
	wire signed [31:0] w_sys_tmp7131;
	wire signed [31:0] w_sys_tmp7133;
	wire signed [31:0] w_sys_tmp7134;
	wire        [31:0] w_sys_tmp7135;
	wire signed [31:0] w_sys_tmp7136;
	wire signed [31:0] w_sys_tmp7137;
	wire signed [31:0] w_sys_tmp7139;
	wire signed [31:0] w_sys_tmp7140;
	wire        [31:0] w_sys_tmp7157;
	wire        [31:0] w_sys_tmp7168;
	wire        [31:0] w_sys_tmp7179;
	wire        [31:0] w_sys_tmp7190;
	wire        [31:0] w_sys_tmp7201;
	wire signed [31:0] w_sys_tmp7204;
	wire signed [31:0] w_sys_tmp7205;
	wire               w_sys_tmp7206;
	wire               w_sys_tmp7207;
	wire signed [31:0] w_sys_tmp7208;
	wire signed [31:0] w_sys_tmp7211;
	wire signed [31:0] w_sys_tmp7212;
	wire        [31:0] w_sys_tmp7213;
	wire signed [31:0] w_sys_tmp7214;
	wire signed [31:0] w_sys_tmp7215;
	wire signed [31:0] w_sys_tmp7217;
	wire signed [31:0] w_sys_tmp7218;
	wire        [31:0] w_sys_tmp7219;
	wire signed [31:0] w_sys_tmp7220;
	wire signed [31:0] w_sys_tmp7221;
	wire signed [31:0] w_sys_tmp7223;
	wire signed [31:0] w_sys_tmp7224;
	wire        [31:0] w_sys_tmp7241;
	wire        [31:0] w_sys_tmp7252;
	wire        [31:0] w_sys_tmp7263;
	wire        [31:0] w_sys_tmp7274;
	wire        [31:0] w_sys_tmp7285;
	wire signed [31:0] w_sys_tmp7288;
	wire signed [31:0] w_sys_tmp7289;
	wire               w_sys_tmp7290;
	wire               w_sys_tmp7291;
	wire signed [31:0] w_sys_tmp7292;
	wire signed [31:0] w_sys_tmp7295;
	wire signed [31:0] w_sys_tmp7296;
	wire        [31:0] w_sys_tmp7297;
	wire signed [31:0] w_sys_tmp7298;
	wire signed [31:0] w_sys_tmp7299;
	wire signed [31:0] w_sys_tmp7301;
	wire signed [31:0] w_sys_tmp7302;
	wire        [31:0] w_sys_tmp7303;
	wire signed [31:0] w_sys_tmp7304;
	wire signed [31:0] w_sys_tmp7305;
	wire signed [31:0] w_sys_tmp7307;
	wire signed [31:0] w_sys_tmp7308;
	wire        [31:0] w_sys_tmp7325;
	wire        [31:0] w_sys_tmp7336;
	wire        [31:0] w_sys_tmp7347;
	wire        [31:0] w_sys_tmp7358;
	wire        [31:0] w_sys_tmp7369;
	wire signed [31:0] w_sys_tmp7372;
	wire signed [31:0] w_sys_tmp7373;
	wire               w_sys_tmp7374;
	wire               w_sys_tmp7375;
	wire signed [31:0] w_sys_tmp7376;
	wire signed [31:0] w_sys_tmp7379;
	wire signed [31:0] w_sys_tmp7380;
	wire        [31:0] w_sys_tmp7381;
	wire signed [31:0] w_sys_tmp7382;
	wire signed [31:0] w_sys_tmp7383;
	wire signed [31:0] w_sys_tmp7385;
	wire signed [31:0] w_sys_tmp7386;
	wire        [31:0] w_sys_tmp7387;
	wire signed [31:0] w_sys_tmp7388;
	wire signed [31:0] w_sys_tmp7389;
	wire signed [31:0] w_sys_tmp7391;
	wire signed [31:0] w_sys_tmp7392;
	wire        [31:0] w_sys_tmp7409;
	wire        [31:0] w_sys_tmp7420;
	wire        [31:0] w_sys_tmp7431;
	wire        [31:0] w_sys_tmp7442;
	wire        [31:0] w_sys_tmp7453;
	wire signed [31:0] w_sys_tmp7456;
	wire               w_sys_tmp7457;
	wire               w_sys_tmp7458;
	wire signed [31:0] w_sys_tmp7459;
	wire signed [31:0] w_sys_tmp7462;
	wire signed [31:0] w_sys_tmp7463;
	wire signed [31:0] w_sys_tmp7464;
	wire signed [31:0] w_sys_tmp7465;
	wire        [31:0] w_sys_tmp7466;
	wire signed [31:0] w_sys_tmp7467;
	wire signed [31:0] w_sys_tmp7468;
	wire signed [31:0] w_sys_tmp7472;
	wire signed [31:0] w_sys_tmp7473;
	wire signed [31:0] w_sys_tmp7475;
	wire        [31:0] w_sys_tmp7476;
	wire signed [31:0] w_sys_tmp7477;
	wire signed [31:0] w_sys_tmp7478;
	wire signed [31:0] w_sys_tmp7482;
	wire signed [31:0] w_sys_tmp7483;
	wire signed [31:0] w_sys_tmp7485;
	wire signed [31:0] w_sys_tmp7486;
	wire signed [31:0] w_sys_tmp7487;
	wire signed [31:0] w_sys_tmp7491;
	wire signed [31:0] w_sys_tmp7492;
	wire signed [31:0] w_sys_tmp7494;
	wire signed [31:0] w_sys_tmp7496;
	wire signed [31:0] w_sys_tmp7497;
	wire signed [31:0] w_sys_tmp7501;
	wire signed [31:0] w_sys_tmp7502;
	wire signed [31:0] w_sys_tmp7504;
	wire signed [31:0] w_sys_tmp7505;
	wire signed [31:0] w_sys_tmp7506;
	wire signed [31:0] w_sys_tmp7510;
	wire signed [31:0] w_sys_tmp7511;
	wire signed [31:0] w_sys_tmp7513;
	wire        [31:0] w_sys_tmp7514;
	wire signed [31:0] w_sys_tmp7515;
	wire signed [31:0] w_sys_tmp7516;
	wire signed [31:0] w_sys_tmp7519;
	wire signed [31:0] w_sys_tmp7520;
	wire signed [31:0] w_sys_tmp7521;
	wire signed [31:0] w_sys_tmp7522;
	wire signed [31:0] w_sys_tmp7523;
	wire signed [31:0] w_sys_tmp7524;
	wire signed [31:0] w_sys_tmp7525;
	wire signed [31:0] w_sys_tmp7526;
	wire signed [31:0] w_sys_tmp7527;
	wire signed [31:0] w_sys_tmp7528;
	wire signed [31:0] w_sys_tmp7529;
	wire signed [31:0] w_sys_tmp7530;
	wire signed [31:0] w_sys_tmp7957;
	wire               w_sys_tmp7958;
	wire               w_sys_tmp7959;
	wire signed [31:0] w_sys_tmp7960;
	wire signed [31:0] w_sys_tmp7963;
	wire signed [31:0] w_sys_tmp7964;
	wire signed [31:0] w_sys_tmp7965;
	wire signed [31:0] w_sys_tmp7966;
	wire        [31:0] w_sys_tmp7967;
	wire signed [31:0] w_sys_tmp7968;
	wire signed [31:0] w_sys_tmp7969;
	wire signed [31:0] w_sys_tmp7973;
	wire signed [31:0] w_sys_tmp7974;
	wire signed [31:0] w_sys_tmp7976;
	wire        [31:0] w_sys_tmp7977;
	wire signed [31:0] w_sys_tmp7978;
	wire signed [31:0] w_sys_tmp7979;
	wire signed [31:0] w_sys_tmp7983;
	wire signed [31:0] w_sys_tmp7984;
	wire signed [31:0] w_sys_tmp7986;
	wire signed [31:0] w_sys_tmp7987;
	wire signed [31:0] w_sys_tmp7988;
	wire signed [31:0] w_sys_tmp7992;
	wire signed [31:0] w_sys_tmp7993;
	wire signed [31:0] w_sys_tmp7995;
	wire signed [31:0] w_sys_tmp7997;
	wire signed [31:0] w_sys_tmp7998;
	wire signed [31:0] w_sys_tmp8002;
	wire signed [31:0] w_sys_tmp8003;
	wire signed [31:0] w_sys_tmp8005;
	wire signed [31:0] w_sys_tmp8006;
	wire signed [31:0] w_sys_tmp8007;
	wire signed [31:0] w_sys_tmp8011;
	wire signed [31:0] w_sys_tmp8012;
	wire signed [31:0] w_sys_tmp8014;
	wire        [31:0] w_sys_tmp8015;
	wire signed [31:0] w_sys_tmp8016;
	wire signed [31:0] w_sys_tmp8017;
	wire signed [31:0] w_sys_tmp8020;
	wire signed [31:0] w_sys_tmp8021;
	wire signed [31:0] w_sys_tmp8022;
	wire signed [31:0] w_sys_tmp8023;
	wire signed [31:0] w_sys_tmp8024;
	wire signed [31:0] w_sys_tmp8025;
	wire signed [31:0] w_sys_tmp8026;
	wire signed [31:0] w_sys_tmp8027;
	wire signed [31:0] w_sys_tmp8028;
	wire signed [31:0] w_sys_tmp8029;
	wire signed [31:0] w_sys_tmp8030;
	wire signed [31:0] w_sys_tmp8031;
	wire signed [31:0] w_sys_tmp8458;
	wire               w_sys_tmp8459;
	wire               w_sys_tmp8460;
	wire signed [31:0] w_sys_tmp8461;
	wire signed [31:0] w_sys_tmp8464;
	wire signed [31:0] w_sys_tmp8465;
	wire signed [31:0] w_sys_tmp8466;
	wire signed [31:0] w_sys_tmp8467;
	wire        [31:0] w_sys_tmp8468;
	wire signed [31:0] w_sys_tmp8469;
	wire signed [31:0] w_sys_tmp8470;
	wire signed [31:0] w_sys_tmp8474;
	wire signed [31:0] w_sys_tmp8475;
	wire signed [31:0] w_sys_tmp8477;
	wire        [31:0] w_sys_tmp8478;
	wire signed [31:0] w_sys_tmp8479;
	wire signed [31:0] w_sys_tmp8480;
	wire signed [31:0] w_sys_tmp8484;
	wire signed [31:0] w_sys_tmp8485;
	wire signed [31:0] w_sys_tmp8487;
	wire signed [31:0] w_sys_tmp8488;
	wire signed [31:0] w_sys_tmp8489;
	wire signed [31:0] w_sys_tmp8493;
	wire signed [31:0] w_sys_tmp8494;
	wire signed [31:0] w_sys_tmp8496;
	wire signed [31:0] w_sys_tmp8498;
	wire signed [31:0] w_sys_tmp8499;
	wire signed [31:0] w_sys_tmp8503;
	wire signed [31:0] w_sys_tmp8504;
	wire signed [31:0] w_sys_tmp8506;
	wire signed [31:0] w_sys_tmp8507;
	wire signed [31:0] w_sys_tmp8508;
	wire signed [31:0] w_sys_tmp8512;
	wire signed [31:0] w_sys_tmp8513;
	wire signed [31:0] w_sys_tmp8515;
	wire        [31:0] w_sys_tmp8516;
	wire signed [31:0] w_sys_tmp8517;
	wire signed [31:0] w_sys_tmp8518;
	wire signed [31:0] w_sys_tmp8521;
	wire signed [31:0] w_sys_tmp8522;
	wire signed [31:0] w_sys_tmp8523;
	wire signed [31:0] w_sys_tmp8524;
	wire signed [31:0] w_sys_tmp8525;
	wire signed [31:0] w_sys_tmp8526;
	wire signed [31:0] w_sys_tmp8527;
	wire signed [31:0] w_sys_tmp8528;
	wire signed [31:0] w_sys_tmp8529;
	wire signed [31:0] w_sys_tmp8530;
	wire signed [31:0] w_sys_tmp8531;
	wire signed [31:0] w_sys_tmp8532;
	wire signed [31:0] w_sys_tmp8959;
	wire               w_sys_tmp8960;
	wire               w_sys_tmp8961;
	wire signed [31:0] w_sys_tmp8962;
	wire signed [31:0] w_sys_tmp8965;
	wire signed [31:0] w_sys_tmp8966;
	wire signed [31:0] w_sys_tmp8967;
	wire signed [31:0] w_sys_tmp8968;
	wire        [31:0] w_sys_tmp8969;
	wire signed [31:0] w_sys_tmp8970;
	wire signed [31:0] w_sys_tmp8971;
	wire signed [31:0] w_sys_tmp8975;
	wire signed [31:0] w_sys_tmp8976;
	wire signed [31:0] w_sys_tmp8978;
	wire        [31:0] w_sys_tmp8979;
	wire signed [31:0] w_sys_tmp8980;
	wire signed [31:0] w_sys_tmp8981;
	wire signed [31:0] w_sys_tmp8985;
	wire signed [31:0] w_sys_tmp8986;
	wire signed [31:0] w_sys_tmp8988;
	wire signed [31:0] w_sys_tmp8989;
	wire signed [31:0] w_sys_tmp8990;
	wire signed [31:0] w_sys_tmp8994;
	wire signed [31:0] w_sys_tmp8995;
	wire signed [31:0] w_sys_tmp8997;
	wire signed [31:0] w_sys_tmp8999;
	wire signed [31:0] w_sys_tmp9000;
	wire signed [31:0] w_sys_tmp9004;
	wire signed [31:0] w_sys_tmp9005;
	wire signed [31:0] w_sys_tmp9007;
	wire signed [31:0] w_sys_tmp9008;
	wire signed [31:0] w_sys_tmp9009;
	wire signed [31:0] w_sys_tmp9013;
	wire signed [31:0] w_sys_tmp9014;
	wire signed [31:0] w_sys_tmp9016;
	wire        [31:0] w_sys_tmp9017;
	wire signed [31:0] w_sys_tmp9018;
	wire signed [31:0] w_sys_tmp9019;
	wire signed [31:0] w_sys_tmp9022;
	wire signed [31:0] w_sys_tmp9023;
	wire signed [31:0] w_sys_tmp9024;
	wire signed [31:0] w_sys_tmp9025;
	wire signed [31:0] w_sys_tmp9026;
	wire signed [31:0] w_sys_tmp9027;
	wire signed [31:0] w_sys_tmp9028;
	wire signed [31:0] w_sys_tmp9029;
	wire signed [31:0] w_sys_tmp9030;
	wire signed [31:0] w_sys_tmp9031;
	wire signed [31:0] w_sys_tmp9032;
	wire signed [31:0] w_sys_tmp9033;
	wire signed [31:0] w_sys_tmp9460;
	wire               w_sys_tmp9461;
	wire               w_sys_tmp9462;
	wire signed [31:0] w_sys_tmp9463;
	wire signed [31:0] w_sys_tmp9466;
	wire signed [31:0] w_sys_tmp9467;
	wire signed [31:0] w_sys_tmp9468;
	wire signed [31:0] w_sys_tmp9469;
	wire        [31:0] w_sys_tmp9470;
	wire signed [31:0] w_sys_tmp9471;
	wire signed [31:0] w_sys_tmp9472;
	wire signed [31:0] w_sys_tmp9476;
	wire signed [31:0] w_sys_tmp9477;
	wire signed [31:0] w_sys_tmp9479;
	wire        [31:0] w_sys_tmp9480;
	wire signed [31:0] w_sys_tmp9481;
	wire signed [31:0] w_sys_tmp9482;
	wire signed [31:0] w_sys_tmp9486;
	wire signed [31:0] w_sys_tmp9487;
	wire signed [31:0] w_sys_tmp9489;
	wire signed [31:0] w_sys_tmp9490;
	wire signed [31:0] w_sys_tmp9491;
	wire signed [31:0] w_sys_tmp9495;
	wire signed [31:0] w_sys_tmp9496;
	wire signed [31:0] w_sys_tmp9498;
	wire signed [31:0] w_sys_tmp9500;
	wire signed [31:0] w_sys_tmp9501;
	wire signed [31:0] w_sys_tmp9505;
	wire signed [31:0] w_sys_tmp9506;
	wire signed [31:0] w_sys_tmp9508;
	wire signed [31:0] w_sys_tmp9509;
	wire signed [31:0] w_sys_tmp9510;
	wire signed [31:0] w_sys_tmp9514;
	wire signed [31:0] w_sys_tmp9515;
	wire signed [31:0] w_sys_tmp9517;
	wire        [31:0] w_sys_tmp9518;
	wire signed [31:0] w_sys_tmp9519;
	wire signed [31:0] w_sys_tmp9520;
	wire signed [31:0] w_sys_tmp9523;
	wire signed [31:0] w_sys_tmp9524;
	wire signed [31:0] w_sys_tmp9525;
	wire signed [31:0] w_sys_tmp9526;
	wire signed [31:0] w_sys_tmp9527;
	wire signed [31:0] w_sys_tmp9528;
	wire signed [31:0] w_sys_tmp9529;
	wire signed [31:0] w_sys_tmp9530;
	wire signed [31:0] w_sys_tmp9531;
	wire signed [31:0] w_sys_tmp9532;
	wire signed [31:0] w_sys_tmp9533;
	wire signed [31:0] w_sys_tmp9534;
	wire signed [31:0] w_sys_tmp9961;
	wire               w_sys_tmp9962;
	wire               w_sys_tmp9963;
	wire signed [31:0] w_sys_tmp9964;
	wire signed [31:0] w_sys_tmp9967;
	wire signed [31:0] w_sys_tmp9968;
	wire signed [31:0] w_sys_tmp9969;
	wire signed [31:0] w_sys_tmp9970;
	wire        [31:0] w_sys_tmp9971;
	wire signed [31:0] w_sys_tmp9972;
	wire signed [31:0] w_sys_tmp9973;
	wire signed [31:0] w_sys_tmp9977;
	wire signed [31:0] w_sys_tmp9978;
	wire signed [31:0] w_sys_tmp9980;
	wire        [31:0] w_sys_tmp9981;
	wire signed [31:0] w_sys_tmp9982;
	wire signed [31:0] w_sys_tmp9983;
	wire signed [31:0] w_sys_tmp9987;
	wire signed [31:0] w_sys_tmp9988;
	wire signed [31:0] w_sys_tmp9990;
	wire signed [31:0] w_sys_tmp9991;
	wire signed [31:0] w_sys_tmp9992;
	wire signed [31:0] w_sys_tmp9996;
	wire signed [31:0] w_sys_tmp9997;
	wire signed [31:0] w_sys_tmp9999;
	wire signed [31:0] w_sys_tmp10001;
	wire signed [31:0] w_sys_tmp10002;
	wire signed [31:0] w_sys_tmp10006;
	wire signed [31:0] w_sys_tmp10007;
	wire signed [31:0] w_sys_tmp10009;
	wire signed [31:0] w_sys_tmp10010;
	wire signed [31:0] w_sys_tmp10011;
	wire signed [31:0] w_sys_tmp10015;
	wire signed [31:0] w_sys_tmp10016;
	wire signed [31:0] w_sys_tmp10018;
	wire        [31:0] w_sys_tmp10019;
	wire signed [31:0] w_sys_tmp10020;
	wire signed [31:0] w_sys_tmp10021;
	wire signed [31:0] w_sys_tmp10024;
	wire signed [31:0] w_sys_tmp10025;
	wire signed [31:0] w_sys_tmp10026;
	wire signed [31:0] w_sys_tmp10027;
	wire signed [31:0] w_sys_tmp10028;
	wire signed [31:0] w_sys_tmp10029;
	wire signed [31:0] w_sys_tmp10030;
	wire signed [31:0] w_sys_tmp10031;
	wire signed [31:0] w_sys_tmp10032;
	wire signed [31:0] w_sys_tmp10033;
	wire signed [31:0] w_sys_tmp10034;
	wire signed [31:0] w_sys_tmp10035;
	wire signed [31:0] w_sys_tmp10462;
	wire               w_sys_tmp10463;
	wire               w_sys_tmp10464;
	wire signed [31:0] w_sys_tmp10465;
	wire signed [31:0] w_sys_tmp10468;
	wire signed [31:0] w_sys_tmp10469;
	wire signed [31:0] w_sys_tmp10470;
	wire signed [31:0] w_sys_tmp10471;
	wire        [31:0] w_sys_tmp10472;
	wire signed [31:0] w_sys_tmp10473;
	wire signed [31:0] w_sys_tmp10474;
	wire signed [31:0] w_sys_tmp10478;
	wire signed [31:0] w_sys_tmp10479;
	wire signed [31:0] w_sys_tmp10481;
	wire        [31:0] w_sys_tmp10482;
	wire signed [31:0] w_sys_tmp10483;
	wire signed [31:0] w_sys_tmp10484;
	wire signed [31:0] w_sys_tmp10488;
	wire signed [31:0] w_sys_tmp10489;
	wire signed [31:0] w_sys_tmp10491;
	wire signed [31:0] w_sys_tmp10492;
	wire signed [31:0] w_sys_tmp10493;
	wire signed [31:0] w_sys_tmp10497;
	wire signed [31:0] w_sys_tmp10498;
	wire signed [31:0] w_sys_tmp10500;
	wire signed [31:0] w_sys_tmp10502;
	wire signed [31:0] w_sys_tmp10503;
	wire signed [31:0] w_sys_tmp10507;
	wire signed [31:0] w_sys_tmp10508;
	wire signed [31:0] w_sys_tmp10510;
	wire signed [31:0] w_sys_tmp10511;
	wire signed [31:0] w_sys_tmp10512;
	wire signed [31:0] w_sys_tmp10516;
	wire signed [31:0] w_sys_tmp10517;
	wire signed [31:0] w_sys_tmp10519;
	wire        [31:0] w_sys_tmp10520;
	wire signed [31:0] w_sys_tmp10521;
	wire signed [31:0] w_sys_tmp10522;
	wire signed [31:0] w_sys_tmp10525;
	wire signed [31:0] w_sys_tmp10526;
	wire signed [31:0] w_sys_tmp10527;
	wire signed [31:0] w_sys_tmp10528;
	wire signed [31:0] w_sys_tmp10529;
	wire signed [31:0] w_sys_tmp10530;
	wire signed [31:0] w_sys_tmp10531;
	wire signed [31:0] w_sys_tmp10532;
	wire signed [31:0] w_sys_tmp10533;
	wire signed [31:0] w_sys_tmp10534;
	wire signed [31:0] w_sys_tmp10535;
	wire signed [31:0] w_sys_tmp10536;
	wire signed [31:0] w_sys_tmp10963;
	wire               w_sys_tmp10964;
	wire               w_sys_tmp10965;
	wire signed [31:0] w_sys_tmp10966;
	wire signed [31:0] w_sys_tmp10969;
	wire signed [31:0] w_sys_tmp10970;
	wire signed [31:0] w_sys_tmp10971;
	wire signed [31:0] w_sys_tmp10972;
	wire        [31:0] w_sys_tmp10973;
	wire signed [31:0] w_sys_tmp10974;
	wire signed [31:0] w_sys_tmp10975;
	wire signed [31:0] w_sys_tmp10979;
	wire signed [31:0] w_sys_tmp10980;
	wire signed [31:0] w_sys_tmp10982;
	wire        [31:0] w_sys_tmp10983;
	wire signed [31:0] w_sys_tmp10984;
	wire signed [31:0] w_sys_tmp10985;
	wire signed [31:0] w_sys_tmp10989;
	wire signed [31:0] w_sys_tmp10990;
	wire signed [31:0] w_sys_tmp10992;
	wire signed [31:0] w_sys_tmp10993;
	wire signed [31:0] w_sys_tmp10994;
	wire signed [31:0] w_sys_tmp10998;
	wire signed [31:0] w_sys_tmp10999;
	wire signed [31:0] w_sys_tmp11001;
	wire signed [31:0] w_sys_tmp11003;
	wire signed [31:0] w_sys_tmp11004;
	wire signed [31:0] w_sys_tmp11008;
	wire signed [31:0] w_sys_tmp11009;
	wire signed [31:0] w_sys_tmp11011;
	wire signed [31:0] w_sys_tmp11012;
	wire signed [31:0] w_sys_tmp11013;
	wire signed [31:0] w_sys_tmp11017;
	wire signed [31:0] w_sys_tmp11018;
	wire signed [31:0] w_sys_tmp11020;
	wire        [31:0] w_sys_tmp11021;
	wire signed [31:0] w_sys_tmp11022;
	wire signed [31:0] w_sys_tmp11023;
	wire signed [31:0] w_sys_tmp11026;
	wire signed [31:0] w_sys_tmp11027;
	wire signed [31:0] w_sys_tmp11028;
	wire signed [31:0] w_sys_tmp11029;
	wire signed [31:0] w_sys_tmp11030;
	wire signed [31:0] w_sys_tmp11031;
	wire signed [31:0] w_sys_tmp11032;
	wire signed [31:0] w_sys_tmp11033;
	wire signed [31:0] w_sys_tmp11034;
	wire signed [31:0] w_sys_tmp11035;
	wire signed [31:0] w_sys_tmp11036;
	wire signed [31:0] w_sys_tmp11037;
	wire signed [31:0] w_sys_tmp11452;
	wire               w_sys_tmp11453;
	wire               w_sys_tmp11454;
	wire signed [31:0] w_sys_tmp11455;
	wire signed [31:0] w_sys_tmp11456;
	wire signed [31:0] w_sys_tmp11457;
	wire               w_sys_tmp11458;
	wire               w_sys_tmp11459;
	wire signed [31:0] w_sys_tmp11460;
	wire signed [31:0] w_sys_tmp11463;
	wire signed [31:0] w_sys_tmp11464;
	wire signed [31:0] w_sys_tmp11465;
	wire        [31:0] w_sys_tmp11466;
	wire signed [31:0] w_sys_tmp11467;
	wire signed [31:0] w_sys_tmp11468;
	wire signed [31:0] w_sys_tmp11470;
	wire signed [31:0] w_sys_tmp11471;
	wire signed [31:0] w_sys_tmp11532;
	wire               w_sys_tmp11533;
	wire               w_sys_tmp11534;
	wire signed [31:0] w_sys_tmp11535;
	wire signed [31:0] w_sys_tmp11537;
	wire signed [31:0] w_sys_tmp11538;
	wire signed [31:0] w_sys_tmp11540;
	wire signed [31:0] w_sys_tmp11541;
	wire signed [31:0] w_sys_tmp11542;
	wire        [31:0] w_sys_tmp11543;
	wire signed [31:0] w_sys_tmp11544;
	wire signed [31:0] w_sys_tmp11545;
	wire signed [31:0] w_sys_tmp11547;
	wire signed [31:0] w_sys_tmp11548;
	wire signed [31:0] w_sys_tmp11549;
	wire signed [31:0] w_sys_tmp11628;
	wire               w_sys_tmp11629;
	wire               w_sys_tmp11630;
	wire signed [31:0] w_sys_tmp11631;
	wire signed [31:0] w_sys_tmp11633;
	wire signed [31:0] w_sys_tmp11634;
	wire signed [31:0] w_sys_tmp11636;
	wire signed [31:0] w_sys_tmp11637;
	wire signed [31:0] w_sys_tmp11638;
	wire        [31:0] w_sys_tmp11639;
	wire signed [31:0] w_sys_tmp11640;
	wire signed [31:0] w_sys_tmp11641;
	wire signed [31:0] w_sys_tmp11643;
	wire signed [31:0] w_sys_tmp11644;
	wire signed [31:0] w_sys_tmp11645;
	wire signed [31:0] w_sys_tmp11724;
	wire               w_sys_tmp11725;
	wire               w_sys_tmp11726;
	wire signed [31:0] w_sys_tmp11727;
	wire signed [31:0] w_sys_tmp11729;
	wire signed [31:0] w_sys_tmp11730;
	wire signed [31:0] w_sys_tmp11732;
	wire signed [31:0] w_sys_tmp11733;
	wire signed [31:0] w_sys_tmp11734;
	wire        [31:0] w_sys_tmp11735;
	wire signed [31:0] w_sys_tmp11736;
	wire signed [31:0] w_sys_tmp11737;
	wire signed [31:0] w_sys_tmp11739;
	wire signed [31:0] w_sys_tmp11740;
	wire signed [31:0] w_sys_tmp11741;
	wire signed [31:0] w_sys_tmp11820;
	wire               w_sys_tmp11821;
	wire               w_sys_tmp11822;
	wire signed [31:0] w_sys_tmp11823;
	wire signed [31:0] w_sys_tmp11825;
	wire signed [31:0] w_sys_tmp11826;
	wire signed [31:0] w_sys_tmp11828;
	wire signed [31:0] w_sys_tmp11829;
	wire signed [31:0] w_sys_tmp11830;
	wire        [31:0] w_sys_tmp11831;
	wire signed [31:0] w_sys_tmp11832;
	wire signed [31:0] w_sys_tmp11833;
	wire signed [31:0] w_sys_tmp11835;
	wire signed [31:0] w_sys_tmp11836;
	wire signed [31:0] w_sys_tmp11837;
	wire signed [31:0] w_sys_tmp11916;
	wire               w_sys_tmp11917;
	wire               w_sys_tmp11918;
	wire signed [31:0] w_sys_tmp11919;
	wire signed [31:0] w_sys_tmp11921;
	wire signed [31:0] w_sys_tmp11922;
	wire signed [31:0] w_sys_tmp11924;
	wire signed [31:0] w_sys_tmp11925;
	wire signed [31:0] w_sys_tmp11926;
	wire        [31:0] w_sys_tmp11927;
	wire signed [31:0] w_sys_tmp11928;
	wire signed [31:0] w_sys_tmp11929;
	wire signed [31:0] w_sys_tmp11931;
	wire signed [31:0] w_sys_tmp11932;
	wire signed [31:0] w_sys_tmp11933;
	wire signed [31:0] w_sys_tmp12012;
	wire               w_sys_tmp12013;
	wire               w_sys_tmp12014;
	wire signed [31:0] w_sys_tmp12015;
	wire signed [31:0] w_sys_tmp12017;
	wire signed [31:0] w_sys_tmp12018;
	wire signed [31:0] w_sys_tmp12020;
	wire signed [31:0] w_sys_tmp12021;
	wire signed [31:0] w_sys_tmp12022;
	wire        [31:0] w_sys_tmp12023;
	wire signed [31:0] w_sys_tmp12024;
	wire signed [31:0] w_sys_tmp12025;
	wire signed [31:0] w_sys_tmp12027;
	wire signed [31:0] w_sys_tmp12028;
	wire signed [31:0] w_sys_tmp12029;
	wire signed [31:0] w_sys_tmp12108;
	wire               w_sys_tmp12109;
	wire               w_sys_tmp12110;
	wire signed [31:0] w_sys_tmp12111;
	wire signed [31:0] w_sys_tmp12113;
	wire signed [31:0] w_sys_tmp12114;
	wire signed [31:0] w_sys_tmp12116;
	wire signed [31:0] w_sys_tmp12117;
	wire signed [31:0] w_sys_tmp12118;
	wire        [31:0] w_sys_tmp12119;
	wire signed [31:0] w_sys_tmp12120;
	wire signed [31:0] w_sys_tmp12121;
	wire signed [31:0] w_sys_tmp12123;
	wire signed [31:0] w_sys_tmp12124;
	wire signed [31:0] w_sys_tmp12125;
	wire signed [31:0] w_sys_tmp12204;
	wire               w_sys_tmp12205;
	wire               w_sys_tmp12206;
	wire signed [31:0] w_sys_tmp12207;
	wire signed [31:0] w_sys_tmp12208;
	wire signed [31:0] w_sys_tmp12209;
	wire               w_sys_tmp12210;
	wire               w_sys_tmp12211;
	wire signed [31:0] w_sys_tmp12212;
	wire signed [31:0] w_sys_tmp12215;
	wire signed [31:0] w_sys_tmp12216;
	wire signed [31:0] w_sys_tmp12217;
	wire        [31:0] w_sys_tmp12218;
	wire signed [31:0] w_sys_tmp12219;
	wire signed [31:0] w_sys_tmp12220;
	wire signed [31:0] w_sys_tmp12222;
	wire signed [31:0] w_sys_tmp12223;
	wire signed [31:0] w_sys_tmp12284;
	wire               w_sys_tmp12285;
	wire               w_sys_tmp12286;
	wire signed [31:0] w_sys_tmp12287;
	wire signed [31:0] w_sys_tmp12289;
	wire signed [31:0] w_sys_tmp12290;
	wire signed [31:0] w_sys_tmp12292;
	wire signed [31:0] w_sys_tmp12293;
	wire signed [31:0] w_sys_tmp12294;
	wire        [31:0] w_sys_tmp12295;
	wire signed [31:0] w_sys_tmp12296;
	wire signed [31:0] w_sys_tmp12297;
	wire signed [31:0] w_sys_tmp12299;
	wire signed [31:0] w_sys_tmp12300;
	wire signed [31:0] w_sys_tmp12301;
	wire signed [31:0] w_sys_tmp12380;
	wire               w_sys_tmp12381;
	wire               w_sys_tmp12382;
	wire signed [31:0] w_sys_tmp12383;
	wire signed [31:0] w_sys_tmp12385;
	wire signed [31:0] w_sys_tmp12386;
	wire signed [31:0] w_sys_tmp12388;
	wire signed [31:0] w_sys_tmp12389;
	wire signed [31:0] w_sys_tmp12390;
	wire        [31:0] w_sys_tmp12391;
	wire signed [31:0] w_sys_tmp12392;
	wire signed [31:0] w_sys_tmp12393;
	wire signed [31:0] w_sys_tmp12395;
	wire signed [31:0] w_sys_tmp12396;
	wire signed [31:0] w_sys_tmp12397;
	wire signed [31:0] w_sys_tmp12476;
	wire               w_sys_tmp12477;
	wire               w_sys_tmp12478;
	wire signed [31:0] w_sys_tmp12479;
	wire signed [31:0] w_sys_tmp12481;
	wire signed [31:0] w_sys_tmp12482;
	wire signed [31:0] w_sys_tmp12484;
	wire signed [31:0] w_sys_tmp12485;
	wire signed [31:0] w_sys_tmp12486;
	wire        [31:0] w_sys_tmp12487;
	wire signed [31:0] w_sys_tmp12488;
	wire signed [31:0] w_sys_tmp12489;
	wire signed [31:0] w_sys_tmp12491;
	wire signed [31:0] w_sys_tmp12492;
	wire signed [31:0] w_sys_tmp12493;
	wire signed [31:0] w_sys_tmp12572;
	wire               w_sys_tmp12573;
	wire               w_sys_tmp12574;
	wire signed [31:0] w_sys_tmp12575;
	wire signed [31:0] w_sys_tmp12577;
	wire signed [31:0] w_sys_tmp12578;
	wire signed [31:0] w_sys_tmp12580;
	wire signed [31:0] w_sys_tmp12581;
	wire signed [31:0] w_sys_tmp12582;
	wire        [31:0] w_sys_tmp12583;
	wire signed [31:0] w_sys_tmp12584;
	wire signed [31:0] w_sys_tmp12585;
	wire signed [31:0] w_sys_tmp12587;
	wire signed [31:0] w_sys_tmp12588;
	wire signed [31:0] w_sys_tmp12589;
	wire signed [31:0] w_sys_tmp12668;
	wire               w_sys_tmp12669;
	wire               w_sys_tmp12670;
	wire signed [31:0] w_sys_tmp12671;
	wire signed [31:0] w_sys_tmp12673;
	wire signed [31:0] w_sys_tmp12674;
	wire signed [31:0] w_sys_tmp12676;
	wire signed [31:0] w_sys_tmp12677;
	wire signed [31:0] w_sys_tmp12678;
	wire        [31:0] w_sys_tmp12679;
	wire signed [31:0] w_sys_tmp12680;
	wire signed [31:0] w_sys_tmp12681;
	wire signed [31:0] w_sys_tmp12683;
	wire signed [31:0] w_sys_tmp12684;
	wire signed [31:0] w_sys_tmp12685;
	wire signed [31:0] w_sys_tmp12764;
	wire               w_sys_tmp12765;
	wire               w_sys_tmp12766;
	wire signed [31:0] w_sys_tmp12767;
	wire signed [31:0] w_sys_tmp12769;
	wire signed [31:0] w_sys_tmp12770;
	wire signed [31:0] w_sys_tmp12772;
	wire signed [31:0] w_sys_tmp12773;
	wire signed [31:0] w_sys_tmp12774;
	wire        [31:0] w_sys_tmp12775;
	wire signed [31:0] w_sys_tmp12776;
	wire signed [31:0] w_sys_tmp12777;
	wire signed [31:0] w_sys_tmp12779;
	wire signed [31:0] w_sys_tmp12780;
	wire signed [31:0] w_sys_tmp12781;
	wire signed [31:0] w_sys_tmp12860;
	wire               w_sys_tmp12861;
	wire               w_sys_tmp12862;
	wire signed [31:0] w_sys_tmp12863;
	wire signed [31:0] w_sys_tmp12865;
	wire signed [31:0] w_sys_tmp12866;
	wire signed [31:0] w_sys_tmp12868;
	wire signed [31:0] w_sys_tmp12869;
	wire signed [31:0] w_sys_tmp12870;
	wire        [31:0] w_sys_tmp12871;
	wire signed [31:0] w_sys_tmp12872;
	wire signed [31:0] w_sys_tmp12873;
	wire signed [31:0] w_sys_tmp12875;
	wire signed [31:0] w_sys_tmp12876;
	wire signed [31:0] w_sys_tmp12877;
	wire signed [31:0] w_sys_tmp12956;
	wire               w_sys_tmp12957;
	wire               w_sys_tmp12958;
	wire signed [31:0] w_sys_tmp12959;
	wire signed [31:0] w_sys_tmp12960;
	wire signed [31:0] w_sys_tmp12961;
	wire               w_sys_tmp12962;
	wire               w_sys_tmp12963;
	wire signed [31:0] w_sys_tmp12964;
	wire signed [31:0] w_sys_tmp12967;
	wire signed [31:0] w_sys_tmp12968;
	wire signed [31:0] w_sys_tmp12969;
	wire        [31:0] w_sys_tmp12970;
	wire signed [31:0] w_sys_tmp12971;
	wire signed [31:0] w_sys_tmp12972;
	wire signed [31:0] w_sys_tmp12974;
	wire signed [31:0] w_sys_tmp12975;
	wire signed [31:0] w_sys_tmp13036;
	wire               w_sys_tmp13037;
	wire               w_sys_tmp13038;
	wire signed [31:0] w_sys_tmp13039;
	wire signed [31:0] w_sys_tmp13041;
	wire signed [31:0] w_sys_tmp13042;
	wire signed [31:0] w_sys_tmp13044;
	wire signed [31:0] w_sys_tmp13045;
	wire signed [31:0] w_sys_tmp13046;
	wire        [31:0] w_sys_tmp13047;
	wire signed [31:0] w_sys_tmp13048;
	wire signed [31:0] w_sys_tmp13049;
	wire signed [31:0] w_sys_tmp13051;
	wire signed [31:0] w_sys_tmp13052;
	wire signed [31:0] w_sys_tmp13053;
	wire signed [31:0] w_sys_tmp13132;
	wire               w_sys_tmp13133;
	wire               w_sys_tmp13134;
	wire signed [31:0] w_sys_tmp13135;
	wire signed [31:0] w_sys_tmp13137;
	wire signed [31:0] w_sys_tmp13138;
	wire signed [31:0] w_sys_tmp13140;
	wire signed [31:0] w_sys_tmp13141;
	wire signed [31:0] w_sys_tmp13142;
	wire        [31:0] w_sys_tmp13143;
	wire signed [31:0] w_sys_tmp13144;
	wire signed [31:0] w_sys_tmp13145;
	wire signed [31:0] w_sys_tmp13147;
	wire signed [31:0] w_sys_tmp13148;
	wire signed [31:0] w_sys_tmp13149;
	wire signed [31:0] w_sys_tmp13228;
	wire               w_sys_tmp13229;
	wire               w_sys_tmp13230;
	wire signed [31:0] w_sys_tmp13231;
	wire signed [31:0] w_sys_tmp13233;
	wire signed [31:0] w_sys_tmp13234;
	wire signed [31:0] w_sys_tmp13236;
	wire signed [31:0] w_sys_tmp13237;
	wire signed [31:0] w_sys_tmp13238;
	wire        [31:0] w_sys_tmp13239;
	wire signed [31:0] w_sys_tmp13240;
	wire signed [31:0] w_sys_tmp13241;
	wire signed [31:0] w_sys_tmp13243;
	wire signed [31:0] w_sys_tmp13244;
	wire signed [31:0] w_sys_tmp13245;
	wire signed [31:0] w_sys_tmp13324;
	wire               w_sys_tmp13325;
	wire               w_sys_tmp13326;
	wire signed [31:0] w_sys_tmp13327;
	wire signed [31:0] w_sys_tmp13329;
	wire signed [31:0] w_sys_tmp13330;
	wire signed [31:0] w_sys_tmp13332;
	wire signed [31:0] w_sys_tmp13333;
	wire signed [31:0] w_sys_tmp13334;
	wire        [31:0] w_sys_tmp13335;
	wire signed [31:0] w_sys_tmp13336;
	wire signed [31:0] w_sys_tmp13337;
	wire signed [31:0] w_sys_tmp13339;
	wire signed [31:0] w_sys_tmp13340;
	wire signed [31:0] w_sys_tmp13341;
	wire signed [31:0] w_sys_tmp13420;
	wire               w_sys_tmp13421;
	wire               w_sys_tmp13422;
	wire signed [31:0] w_sys_tmp13423;
	wire signed [31:0] w_sys_tmp13425;
	wire signed [31:0] w_sys_tmp13426;
	wire signed [31:0] w_sys_tmp13428;
	wire signed [31:0] w_sys_tmp13429;
	wire signed [31:0] w_sys_tmp13430;
	wire        [31:0] w_sys_tmp13431;
	wire signed [31:0] w_sys_tmp13432;
	wire signed [31:0] w_sys_tmp13433;
	wire signed [31:0] w_sys_tmp13435;
	wire signed [31:0] w_sys_tmp13436;
	wire signed [31:0] w_sys_tmp13437;
	wire signed [31:0] w_sys_tmp13516;
	wire               w_sys_tmp13517;
	wire               w_sys_tmp13518;
	wire signed [31:0] w_sys_tmp13519;
	wire signed [31:0] w_sys_tmp13521;
	wire signed [31:0] w_sys_tmp13522;
	wire signed [31:0] w_sys_tmp13524;
	wire signed [31:0] w_sys_tmp13525;
	wire signed [31:0] w_sys_tmp13526;
	wire        [31:0] w_sys_tmp13527;
	wire signed [31:0] w_sys_tmp13528;
	wire signed [31:0] w_sys_tmp13529;
	wire signed [31:0] w_sys_tmp13531;
	wire signed [31:0] w_sys_tmp13532;
	wire signed [31:0] w_sys_tmp13533;
	wire signed [31:0] w_sys_tmp13612;
	wire               w_sys_tmp13613;
	wire               w_sys_tmp13614;
	wire signed [31:0] w_sys_tmp13615;
	wire signed [31:0] w_sys_tmp13617;
	wire signed [31:0] w_sys_tmp13618;
	wire signed [31:0] w_sys_tmp13620;
	wire signed [31:0] w_sys_tmp13621;
	wire signed [31:0] w_sys_tmp13622;
	wire        [31:0] w_sys_tmp13623;
	wire signed [31:0] w_sys_tmp13624;
	wire signed [31:0] w_sys_tmp13625;
	wire signed [31:0] w_sys_tmp13627;
	wire signed [31:0] w_sys_tmp13628;
	wire signed [31:0] w_sys_tmp13629;
	wire signed [31:0] w_sys_tmp13708;
	wire               w_sys_tmp13709;
	wire               w_sys_tmp13710;
	wire signed [31:0] w_sys_tmp13711;
	wire signed [31:0] w_sys_tmp13712;
	wire signed [31:0] w_sys_tmp13713;
	wire               w_sys_tmp13714;
	wire               w_sys_tmp13715;
	wire signed [31:0] w_sys_tmp13716;
	wire signed [31:0] w_sys_tmp13719;
	wire signed [31:0] w_sys_tmp13720;
	wire signed [31:0] w_sys_tmp13721;
	wire        [31:0] w_sys_tmp13722;
	wire signed [31:0] w_sys_tmp13723;
	wire signed [31:0] w_sys_tmp13724;
	wire signed [31:0] w_sys_tmp13726;
	wire signed [31:0] w_sys_tmp13727;
	wire signed [31:0] w_sys_tmp13788;
	wire               w_sys_tmp13789;
	wire               w_sys_tmp13790;
	wire signed [31:0] w_sys_tmp13791;
	wire signed [31:0] w_sys_tmp13793;
	wire signed [31:0] w_sys_tmp13794;
	wire signed [31:0] w_sys_tmp13796;
	wire signed [31:0] w_sys_tmp13797;
	wire signed [31:0] w_sys_tmp13798;
	wire        [31:0] w_sys_tmp13799;
	wire signed [31:0] w_sys_tmp13800;
	wire signed [31:0] w_sys_tmp13801;
	wire signed [31:0] w_sys_tmp13803;
	wire signed [31:0] w_sys_tmp13804;
	wire signed [31:0] w_sys_tmp13805;
	wire signed [31:0] w_sys_tmp13884;
	wire               w_sys_tmp13885;
	wire               w_sys_tmp13886;
	wire signed [31:0] w_sys_tmp13887;
	wire signed [31:0] w_sys_tmp13889;
	wire signed [31:0] w_sys_tmp13890;
	wire signed [31:0] w_sys_tmp13892;
	wire signed [31:0] w_sys_tmp13893;
	wire signed [31:0] w_sys_tmp13894;
	wire        [31:0] w_sys_tmp13895;
	wire signed [31:0] w_sys_tmp13896;
	wire signed [31:0] w_sys_tmp13897;
	wire signed [31:0] w_sys_tmp13899;
	wire signed [31:0] w_sys_tmp13900;
	wire signed [31:0] w_sys_tmp13901;
	wire signed [31:0] w_sys_tmp13980;
	wire               w_sys_tmp13981;
	wire               w_sys_tmp13982;
	wire signed [31:0] w_sys_tmp13983;
	wire signed [31:0] w_sys_tmp13985;
	wire signed [31:0] w_sys_tmp13986;
	wire signed [31:0] w_sys_tmp13988;
	wire signed [31:0] w_sys_tmp13989;
	wire signed [31:0] w_sys_tmp13990;
	wire        [31:0] w_sys_tmp13991;
	wire signed [31:0] w_sys_tmp13992;
	wire signed [31:0] w_sys_tmp13993;
	wire signed [31:0] w_sys_tmp13995;
	wire signed [31:0] w_sys_tmp13996;
	wire signed [31:0] w_sys_tmp13997;
	wire signed [31:0] w_sys_tmp14076;
	wire               w_sys_tmp14077;
	wire               w_sys_tmp14078;
	wire signed [31:0] w_sys_tmp14079;
	wire signed [31:0] w_sys_tmp14081;
	wire signed [31:0] w_sys_tmp14082;
	wire signed [31:0] w_sys_tmp14084;
	wire signed [31:0] w_sys_tmp14085;
	wire signed [31:0] w_sys_tmp14086;
	wire        [31:0] w_sys_tmp14087;
	wire signed [31:0] w_sys_tmp14088;
	wire signed [31:0] w_sys_tmp14089;
	wire signed [31:0] w_sys_tmp14091;
	wire signed [31:0] w_sys_tmp14092;
	wire signed [31:0] w_sys_tmp14093;
	wire signed [31:0] w_sys_tmp14172;
	wire               w_sys_tmp14173;
	wire               w_sys_tmp14174;
	wire signed [31:0] w_sys_tmp14175;
	wire signed [31:0] w_sys_tmp14177;
	wire signed [31:0] w_sys_tmp14178;
	wire signed [31:0] w_sys_tmp14180;
	wire signed [31:0] w_sys_tmp14181;
	wire signed [31:0] w_sys_tmp14182;
	wire        [31:0] w_sys_tmp14183;
	wire signed [31:0] w_sys_tmp14184;
	wire signed [31:0] w_sys_tmp14185;
	wire signed [31:0] w_sys_tmp14187;
	wire signed [31:0] w_sys_tmp14188;
	wire signed [31:0] w_sys_tmp14189;
	wire signed [31:0] w_sys_tmp14268;
	wire               w_sys_tmp14269;
	wire               w_sys_tmp14270;
	wire signed [31:0] w_sys_tmp14271;
	wire signed [31:0] w_sys_tmp14273;
	wire signed [31:0] w_sys_tmp14274;
	wire signed [31:0] w_sys_tmp14276;
	wire signed [31:0] w_sys_tmp14277;
	wire signed [31:0] w_sys_tmp14278;
	wire        [31:0] w_sys_tmp14279;
	wire signed [31:0] w_sys_tmp14280;
	wire signed [31:0] w_sys_tmp14281;
	wire signed [31:0] w_sys_tmp14283;
	wire signed [31:0] w_sys_tmp14284;
	wire signed [31:0] w_sys_tmp14285;
	wire signed [31:0] w_sys_tmp14364;
	wire               w_sys_tmp14365;
	wire               w_sys_tmp14366;
	wire signed [31:0] w_sys_tmp14367;
	wire signed [31:0] w_sys_tmp14369;
	wire signed [31:0] w_sys_tmp14370;
	wire signed [31:0] w_sys_tmp14372;
	wire signed [31:0] w_sys_tmp14373;
	wire signed [31:0] w_sys_tmp14374;
	wire        [31:0] w_sys_tmp14375;
	wire signed [31:0] w_sys_tmp14376;
	wire signed [31:0] w_sys_tmp14377;
	wire signed [31:0] w_sys_tmp14379;
	wire signed [31:0] w_sys_tmp14380;
	wire signed [31:0] w_sys_tmp14381;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 6'h1);
	assign w_fld_T_0_addr_0 = 15'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 15'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 15'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_fld_V_3_addr_0 = 15'sh0;
	assign w_fld_V_3_datain_0 = 32'h0;
	assign w_fld_V_3_r_w_0 = 1'h0;
	assign w_fld_V_3_ce_0 = w_sys_ce;
	assign w_fld_V_3_ce_1 = w_sys_ce;
	assign w_sub19_T_addr = ( (|r_sys_processing_methodID) ? r_sub19_T_addr : 15'sh0 ) ;
	assign w_sub19_T_datain = ( (|r_sys_processing_methodID) ? r_sub19_T_datain : 32'h0 ) ;
	assign w_sub19_T_r_w = ( (|r_sys_processing_methodID) ? r_sub19_T_r_w : 1'h0 ) ;
	assign w_sub19_V_addr = ( (|r_sys_processing_methodID) ? r_sub19_V_addr : 15'sh0 ) ;
	assign w_sub19_V_datain = ( (|r_sys_processing_methodID) ? r_sub19_V_datain : 32'h0 ) ;
	assign w_sub19_V_r_w = ( (|r_sys_processing_methodID) ? r_sub19_V_r_w : 1'h0 ) ;
	assign w_sub19_U_addr = ( (|r_sys_processing_methodID) ? r_sub19_U_addr : 15'sh0 ) ;
	assign w_sub19_U_datain = ( (|r_sys_processing_methodID) ? r_sub19_U_datain : 32'h0 ) ;
	assign w_sub19_U_r_w = ( (|r_sys_processing_methodID) ? r_sub19_U_r_w : 1'h0 ) ;
	assign w_sub19_result_addr = ( (|r_sys_processing_methodID) ? r_sub19_result_addr : 15'sh0 ) ;
	assign w_sub19_result_datain = ( (|r_sys_processing_methodID) ? r_sub19_result_datain : 32'h0 ) ;
	assign w_sub19_result_r_w = ( (|r_sys_processing_methodID) ? r_sub19_result_r_w : 1'h0 ) ;
	assign w_sub12_T_addr = ( (|r_sys_processing_methodID) ? r_sub12_T_addr : 15'sh0 ) ;
	assign w_sub12_T_datain = ( (|r_sys_processing_methodID) ? r_sub12_T_datain : 32'h0 ) ;
	assign w_sub12_T_r_w = ( (|r_sys_processing_methodID) ? r_sub12_T_r_w : 1'h0 ) ;
	assign w_sub12_V_addr = ( (|r_sys_processing_methodID) ? r_sub12_V_addr : 15'sh0 ) ;
	assign w_sub12_V_datain = ( (|r_sys_processing_methodID) ? r_sub12_V_datain : 32'h0 ) ;
	assign w_sub12_V_r_w = ( (|r_sys_processing_methodID) ? r_sub12_V_r_w : 1'h0 ) ;
	assign w_sub12_U_addr = ( (|r_sys_processing_methodID) ? r_sub12_U_addr : 15'sh0 ) ;
	assign w_sub12_U_datain = ( (|r_sys_processing_methodID) ? r_sub12_U_datain : 32'h0 ) ;
	assign w_sub12_U_r_w = ( (|r_sys_processing_methodID) ? r_sub12_U_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 15'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub11_T_addr = ( (|r_sys_processing_methodID) ? r_sub11_T_addr : 15'sh0 ) ;
	assign w_sub11_T_datain = ( (|r_sys_processing_methodID) ? r_sub11_T_datain : 32'h0 ) ;
	assign w_sub11_T_r_w = ( (|r_sys_processing_methodID) ? r_sub11_T_r_w : 1'h0 ) ;
	assign w_sub11_V_addr = ( (|r_sys_processing_methodID) ? r_sub11_V_addr : 15'sh0 ) ;
	assign w_sub11_V_datain = ( (|r_sys_processing_methodID) ? r_sub11_V_datain : 32'h0 ) ;
	assign w_sub11_V_r_w = ( (|r_sys_processing_methodID) ? r_sub11_V_r_w : 1'h0 ) ;
	assign w_sub11_U_addr = ( (|r_sys_processing_methodID) ? r_sub11_U_addr : 15'sh0 ) ;
	assign w_sub11_U_datain = ( (|r_sys_processing_methodID) ? r_sub11_U_datain : 32'h0 ) ;
	assign w_sub11_U_r_w = ( (|r_sys_processing_methodID) ? r_sub11_U_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 15'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_T_addr = ( (|r_sys_processing_methodID) ? r_sub14_T_addr : 15'sh0 ) ;
	assign w_sub14_T_datain = ( (|r_sys_processing_methodID) ? r_sub14_T_datain : 32'h0 ) ;
	assign w_sub14_T_r_w = ( (|r_sys_processing_methodID) ? r_sub14_T_r_w : 1'h0 ) ;
	assign w_sub14_V_addr = ( (|r_sys_processing_methodID) ? r_sub14_V_addr : 15'sh0 ) ;
	assign w_sub14_V_datain = ( (|r_sys_processing_methodID) ? r_sub14_V_datain : 32'h0 ) ;
	assign w_sub14_V_r_w = ( (|r_sys_processing_methodID) ? r_sub14_V_r_w : 1'h0 ) ;
	assign w_sub14_U_addr = ( (|r_sys_processing_methodID) ? r_sub14_U_addr : 15'sh0 ) ;
	assign w_sub14_U_datain = ( (|r_sys_processing_methodID) ? r_sub14_U_datain : 32'h0 ) ;
	assign w_sub14_U_r_w = ( (|r_sys_processing_methodID) ? r_sub14_U_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 15'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub13_T_addr = ( (|r_sys_processing_methodID) ? r_sub13_T_addr : 15'sh0 ) ;
	assign w_sub13_T_datain = ( (|r_sys_processing_methodID) ? r_sub13_T_datain : 32'h0 ) ;
	assign w_sub13_T_r_w = ( (|r_sys_processing_methodID) ? r_sub13_T_r_w : 1'h0 ) ;
	assign w_sub13_V_addr = ( (|r_sys_processing_methodID) ? r_sub13_V_addr : 15'sh0 ) ;
	assign w_sub13_V_datain = ( (|r_sys_processing_methodID) ? r_sub13_V_datain : 32'h0 ) ;
	assign w_sub13_V_r_w = ( (|r_sys_processing_methodID) ? r_sub13_V_r_w : 1'h0 ) ;
	assign w_sub13_U_addr = ( (|r_sys_processing_methodID) ? r_sub13_U_addr : 15'sh0 ) ;
	assign w_sub13_U_datain = ( (|r_sys_processing_methodID) ? r_sub13_U_datain : 32'h0 ) ;
	assign w_sub13_U_r_w = ( (|r_sys_processing_methodID) ? r_sub13_U_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 15'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub16_T_addr = ( (|r_sys_processing_methodID) ? r_sub16_T_addr : 15'sh0 ) ;
	assign w_sub16_T_datain = ( (|r_sys_processing_methodID) ? r_sub16_T_datain : 32'h0 ) ;
	assign w_sub16_T_r_w = ( (|r_sys_processing_methodID) ? r_sub16_T_r_w : 1'h0 ) ;
	assign w_sub16_V_addr = ( (|r_sys_processing_methodID) ? r_sub16_V_addr : 15'sh0 ) ;
	assign w_sub16_V_datain = ( (|r_sys_processing_methodID) ? r_sub16_V_datain : 32'h0 ) ;
	assign w_sub16_V_r_w = ( (|r_sys_processing_methodID) ? r_sub16_V_r_w : 1'h0 ) ;
	assign w_sub16_U_addr = ( (|r_sys_processing_methodID) ? r_sub16_U_addr : 15'sh0 ) ;
	assign w_sub16_U_datain = ( (|r_sys_processing_methodID) ? r_sub16_U_datain : 32'h0 ) ;
	assign w_sub16_U_r_w = ( (|r_sys_processing_methodID) ? r_sub16_U_r_w : 1'h0 ) ;
	assign w_sub16_result_addr = ( (|r_sys_processing_methodID) ? r_sub16_result_addr : 15'sh0 ) ;
	assign w_sub16_result_datain = ( (|r_sys_processing_methodID) ? r_sub16_result_datain : 32'h0 ) ;
	assign w_sub16_result_r_w = ( (|r_sys_processing_methodID) ? r_sub16_result_r_w : 1'h0 ) ;
	assign w_sub15_T_addr = ( (|r_sys_processing_methodID) ? r_sub15_T_addr : 15'sh0 ) ;
	assign w_sub15_T_datain = ( (|r_sys_processing_methodID) ? r_sub15_T_datain : 32'h0 ) ;
	assign w_sub15_T_r_w = ( (|r_sys_processing_methodID) ? r_sub15_T_r_w : 1'h0 ) ;
	assign w_sub15_V_addr = ( (|r_sys_processing_methodID) ? r_sub15_V_addr : 15'sh0 ) ;
	assign w_sub15_V_datain = ( (|r_sys_processing_methodID) ? r_sub15_V_datain : 32'h0 ) ;
	assign w_sub15_V_r_w = ( (|r_sys_processing_methodID) ? r_sub15_V_r_w : 1'h0 ) ;
	assign w_sub15_U_addr = ( (|r_sys_processing_methodID) ? r_sub15_U_addr : 15'sh0 ) ;
	assign w_sub15_U_datain = ( (|r_sys_processing_methodID) ? r_sub15_U_datain : 32'h0 ) ;
	assign w_sub15_U_r_w = ( (|r_sys_processing_methodID) ? r_sub15_U_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 15'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub18_T_addr = ( (|r_sys_processing_methodID) ? r_sub18_T_addr : 15'sh0 ) ;
	assign w_sub18_T_datain = ( (|r_sys_processing_methodID) ? r_sub18_T_datain : 32'h0 ) ;
	assign w_sub18_T_r_w = ( (|r_sys_processing_methodID) ? r_sub18_T_r_w : 1'h0 ) ;
	assign w_sub18_V_addr = ( (|r_sys_processing_methodID) ? r_sub18_V_addr : 15'sh0 ) ;
	assign w_sub18_V_datain = ( (|r_sys_processing_methodID) ? r_sub18_V_datain : 32'h0 ) ;
	assign w_sub18_V_r_w = ( (|r_sys_processing_methodID) ? r_sub18_V_r_w : 1'h0 ) ;
	assign w_sub18_U_addr = ( (|r_sys_processing_methodID) ? r_sub18_U_addr : 15'sh0 ) ;
	assign w_sub18_U_datain = ( (|r_sys_processing_methodID) ? r_sub18_U_datain : 32'h0 ) ;
	assign w_sub18_U_r_w = ( (|r_sys_processing_methodID) ? r_sub18_U_r_w : 1'h0 ) ;
	assign w_sub18_result_addr = ( (|r_sys_processing_methodID) ? r_sub18_result_addr : 15'sh0 ) ;
	assign w_sub18_result_datain = ( (|r_sys_processing_methodID) ? r_sub18_result_datain : 32'h0 ) ;
	assign w_sub18_result_r_w = ( (|r_sys_processing_methodID) ? r_sub18_result_r_w : 1'h0 ) ;
	assign w_sub17_T_addr = ( (|r_sys_processing_methodID) ? r_sub17_T_addr : 15'sh0 ) ;
	assign w_sub17_T_datain = ( (|r_sys_processing_methodID) ? r_sub17_T_datain : 32'h0 ) ;
	assign w_sub17_T_r_w = ( (|r_sys_processing_methodID) ? r_sub17_T_r_w : 1'h0 ) ;
	assign w_sub17_V_addr = ( (|r_sys_processing_methodID) ? r_sub17_V_addr : 15'sh0 ) ;
	assign w_sub17_V_datain = ( (|r_sys_processing_methodID) ? r_sub17_V_datain : 32'h0 ) ;
	assign w_sub17_V_r_w = ( (|r_sys_processing_methodID) ? r_sub17_V_r_w : 1'h0 ) ;
	assign w_sub17_U_addr = ( (|r_sys_processing_methodID) ? r_sub17_U_addr : 15'sh0 ) ;
	assign w_sub17_U_datain = ( (|r_sys_processing_methodID) ? r_sub17_U_datain : 32'h0 ) ;
	assign w_sub17_U_r_w = ( (|r_sys_processing_methodID) ? r_sub17_U_r_w : 1'h0 ) ;
	assign w_sub17_result_addr = ( (|r_sys_processing_methodID) ? r_sub17_result_addr : 15'sh0 ) ;
	assign w_sub17_result_datain = ( (|r_sys_processing_methodID) ? r_sub17_result_datain : 32'h0 ) ;
	assign w_sub17_result_r_w = ( (|r_sys_processing_methodID) ? r_sub17_result_r_w : 1'h0 ) ;
	assign w_sub20_T_addr = ( (|r_sys_processing_methodID) ? r_sub20_T_addr : 15'sh0 ) ;
	assign w_sub20_T_datain = ( (|r_sys_processing_methodID) ? r_sub20_T_datain : 32'h0 ) ;
	assign w_sub20_T_r_w = ( (|r_sys_processing_methodID) ? r_sub20_T_r_w : 1'h0 ) ;
	assign w_sub20_V_addr = ( (|r_sys_processing_methodID) ? r_sub20_V_addr : 15'sh0 ) ;
	assign w_sub20_V_datain = ( (|r_sys_processing_methodID) ? r_sub20_V_datain : 32'h0 ) ;
	assign w_sub20_V_r_w = ( (|r_sys_processing_methodID) ? r_sub20_V_r_w : 1'h0 ) ;
	assign w_sub20_U_addr = ( (|r_sys_processing_methodID) ? r_sub20_U_addr : 15'sh0 ) ;
	assign w_sub20_U_datain = ( (|r_sys_processing_methodID) ? r_sub20_U_datain : 32'h0 ) ;
	assign w_sub20_U_r_w = ( (|r_sys_processing_methodID) ? r_sub20_U_r_w : 1'h0 ) ;
	assign w_sub20_result_addr = ( (|r_sys_processing_methodID) ? r_sub20_result_addr : 15'sh0 ) ;
	assign w_sub20_result_datain = ( (|r_sys_processing_methodID) ? r_sub20_result_datain : 32'h0 ) ;
	assign w_sub20_result_r_w = ( (|r_sys_processing_methodID) ? r_sub20_result_r_w : 1'h0 ) ;
	assign w_sub21_T_addr = ( (|r_sys_processing_methodID) ? r_sub21_T_addr : 15'sh0 ) ;
	assign w_sub21_T_datain = ( (|r_sys_processing_methodID) ? r_sub21_T_datain : 32'h0 ) ;
	assign w_sub21_T_r_w = ( (|r_sys_processing_methodID) ? r_sub21_T_r_w : 1'h0 ) ;
	assign w_sub21_V_addr = ( (|r_sys_processing_methodID) ? r_sub21_V_addr : 15'sh0 ) ;
	assign w_sub21_V_datain = ( (|r_sys_processing_methodID) ? r_sub21_V_datain : 32'h0 ) ;
	assign w_sub21_V_r_w = ( (|r_sys_processing_methodID) ? r_sub21_V_r_w : 1'h0 ) ;
	assign w_sub21_U_addr = ( (|r_sys_processing_methodID) ? r_sub21_U_addr : 15'sh0 ) ;
	assign w_sub21_U_datain = ( (|r_sys_processing_methodID) ? r_sub21_U_datain : 32'h0 ) ;
	assign w_sub21_U_r_w = ( (|r_sys_processing_methodID) ? r_sub21_U_r_w : 1'h0 ) ;
	assign w_sub21_result_addr = ( (|r_sys_processing_methodID) ? r_sub21_result_addr : 15'sh0 ) ;
	assign w_sub21_result_datain = ( (|r_sys_processing_methodID) ? r_sub21_result_datain : 32'h0 ) ;
	assign w_sub21_result_r_w = ( (|r_sys_processing_methodID) ? r_sub21_result_r_w : 1'h0 ) ;
	assign w_sub28_T_addr = ( (|r_sys_processing_methodID) ? r_sub28_T_addr : 15'sh0 ) ;
	assign w_sub28_T_datain = ( (|r_sys_processing_methodID) ? r_sub28_T_datain : 32'h0 ) ;
	assign w_sub28_T_r_w = ( (|r_sys_processing_methodID) ? r_sub28_T_r_w : 1'h0 ) ;
	assign w_sub28_V_addr = ( (|r_sys_processing_methodID) ? r_sub28_V_addr : 15'sh0 ) ;
	assign w_sub28_V_datain = ( (|r_sys_processing_methodID) ? r_sub28_V_datain : 32'h0 ) ;
	assign w_sub28_V_r_w = ( (|r_sys_processing_methodID) ? r_sub28_V_r_w : 1'h0 ) ;
	assign w_sub28_U_addr = ( (|r_sys_processing_methodID) ? r_sub28_U_addr : 15'sh0 ) ;
	assign w_sub28_U_datain = ( (|r_sys_processing_methodID) ? r_sub28_U_datain : 32'h0 ) ;
	assign w_sub28_U_r_w = ( (|r_sys_processing_methodID) ? r_sub28_U_r_w : 1'h0 ) ;
	assign w_sub28_result_addr = ( (|r_sys_processing_methodID) ? r_sub28_result_addr : 15'sh0 ) ;
	assign w_sub28_result_datain = ( (|r_sys_processing_methodID) ? r_sub28_result_datain : 32'h0 ) ;
	assign w_sub28_result_r_w = ( (|r_sys_processing_methodID) ? r_sub28_result_r_w : 1'h0 ) ;
	assign w_sub29_T_addr = ( (|r_sys_processing_methodID) ? r_sub29_T_addr : 15'sh0 ) ;
	assign w_sub29_T_datain = ( (|r_sys_processing_methodID) ? r_sub29_T_datain : 32'h0 ) ;
	assign w_sub29_T_r_w = ( (|r_sys_processing_methodID) ? r_sub29_T_r_w : 1'h0 ) ;
	assign w_sub29_V_addr = ( (|r_sys_processing_methodID) ? r_sub29_V_addr : 15'sh0 ) ;
	assign w_sub29_V_datain = ( (|r_sys_processing_methodID) ? r_sub29_V_datain : 32'h0 ) ;
	assign w_sub29_V_r_w = ( (|r_sys_processing_methodID) ? r_sub29_V_r_w : 1'h0 ) ;
	assign w_sub29_U_addr = ( (|r_sys_processing_methodID) ? r_sub29_U_addr : 15'sh0 ) ;
	assign w_sub29_U_datain = ( (|r_sys_processing_methodID) ? r_sub29_U_datain : 32'h0 ) ;
	assign w_sub29_U_r_w = ( (|r_sys_processing_methodID) ? r_sub29_U_r_w : 1'h0 ) ;
	assign w_sub29_result_addr = ( (|r_sys_processing_methodID) ? r_sub29_result_addr : 15'sh0 ) ;
	assign w_sub29_result_datain = ( (|r_sys_processing_methodID) ? r_sub29_result_datain : 32'h0 ) ;
	assign w_sub29_result_r_w = ( (|r_sys_processing_methodID) ? r_sub29_result_r_w : 1'h0 ) ;
	assign w_sub26_T_addr = ( (|r_sys_processing_methodID) ? r_sub26_T_addr : 15'sh0 ) ;
	assign w_sub26_T_datain = ( (|r_sys_processing_methodID) ? r_sub26_T_datain : 32'h0 ) ;
	assign w_sub26_T_r_w = ( (|r_sys_processing_methodID) ? r_sub26_T_r_w : 1'h0 ) ;
	assign w_sub26_V_addr = ( (|r_sys_processing_methodID) ? r_sub26_V_addr : 15'sh0 ) ;
	assign w_sub26_V_datain = ( (|r_sys_processing_methodID) ? r_sub26_V_datain : 32'h0 ) ;
	assign w_sub26_V_r_w = ( (|r_sys_processing_methodID) ? r_sub26_V_r_w : 1'h0 ) ;
	assign w_sub26_U_addr = ( (|r_sys_processing_methodID) ? r_sub26_U_addr : 15'sh0 ) ;
	assign w_sub26_U_datain = ( (|r_sys_processing_methodID) ? r_sub26_U_datain : 32'h0 ) ;
	assign w_sub26_U_r_w = ( (|r_sys_processing_methodID) ? r_sub26_U_r_w : 1'h0 ) ;
	assign w_sub26_result_addr = ( (|r_sys_processing_methodID) ? r_sub26_result_addr : 15'sh0 ) ;
	assign w_sub26_result_datain = ( (|r_sys_processing_methodID) ? r_sub26_result_datain : 32'h0 ) ;
	assign w_sub26_result_r_w = ( (|r_sys_processing_methodID) ? r_sub26_result_r_w : 1'h0 ) ;
	assign w_sub09_T_addr = ( (|r_sys_processing_methodID) ? r_sub09_T_addr : 15'sh0 ) ;
	assign w_sub09_T_datain = ( (|r_sys_processing_methodID) ? r_sub09_T_datain : 32'h0 ) ;
	assign w_sub09_T_r_w = ( (|r_sys_processing_methodID) ? r_sub09_T_r_w : 1'h0 ) ;
	assign w_sub09_V_addr = ( (|r_sys_processing_methodID) ? r_sub09_V_addr : 15'sh0 ) ;
	assign w_sub09_V_datain = ( (|r_sys_processing_methodID) ? r_sub09_V_datain : 32'h0 ) ;
	assign w_sub09_V_r_w = ( (|r_sys_processing_methodID) ? r_sub09_V_r_w : 1'h0 ) ;
	assign w_sub09_U_addr = ( (|r_sys_processing_methodID) ? r_sub09_U_addr : 15'sh0 ) ;
	assign w_sub09_U_datain = ( (|r_sys_processing_methodID) ? r_sub09_U_datain : 32'h0 ) ;
	assign w_sub09_U_r_w = ( (|r_sys_processing_methodID) ? r_sub09_U_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 15'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub27_T_addr = ( (|r_sys_processing_methodID) ? r_sub27_T_addr : 15'sh0 ) ;
	assign w_sub27_T_datain = ( (|r_sys_processing_methodID) ? r_sub27_T_datain : 32'h0 ) ;
	assign w_sub27_T_r_w = ( (|r_sys_processing_methodID) ? r_sub27_T_r_w : 1'h0 ) ;
	assign w_sub27_V_addr = ( (|r_sys_processing_methodID) ? r_sub27_V_addr : 15'sh0 ) ;
	assign w_sub27_V_datain = ( (|r_sys_processing_methodID) ? r_sub27_V_datain : 32'h0 ) ;
	assign w_sub27_V_r_w = ( (|r_sys_processing_methodID) ? r_sub27_V_r_w : 1'h0 ) ;
	assign w_sub27_U_addr = ( (|r_sys_processing_methodID) ? r_sub27_U_addr : 15'sh0 ) ;
	assign w_sub27_U_datain = ( (|r_sys_processing_methodID) ? r_sub27_U_datain : 32'h0 ) ;
	assign w_sub27_U_r_w = ( (|r_sys_processing_methodID) ? r_sub27_U_r_w : 1'h0 ) ;
	assign w_sub27_result_addr = ( (|r_sys_processing_methodID) ? r_sub27_result_addr : 15'sh0 ) ;
	assign w_sub27_result_datain = ( (|r_sys_processing_methodID) ? r_sub27_result_datain : 32'h0 ) ;
	assign w_sub27_result_r_w = ( (|r_sys_processing_methodID) ? r_sub27_result_r_w : 1'h0 ) ;
	assign w_sub08_T_addr = ( (|r_sys_processing_methodID) ? r_sub08_T_addr : 15'sh0 ) ;
	assign w_sub08_T_datain = ( (|r_sys_processing_methodID) ? r_sub08_T_datain : 32'h0 ) ;
	assign w_sub08_T_r_w = ( (|r_sys_processing_methodID) ? r_sub08_T_r_w : 1'h0 ) ;
	assign w_sub08_V_addr = ( (|r_sys_processing_methodID) ? r_sub08_V_addr : 15'sh0 ) ;
	assign w_sub08_V_datain = ( (|r_sys_processing_methodID) ? r_sub08_V_datain : 32'h0 ) ;
	assign w_sub08_V_r_w = ( (|r_sys_processing_methodID) ? r_sub08_V_r_w : 1'h0 ) ;
	assign w_sub08_U_addr = ( (|r_sys_processing_methodID) ? r_sub08_U_addr : 15'sh0 ) ;
	assign w_sub08_U_datain = ( (|r_sys_processing_methodID) ? r_sub08_U_datain : 32'h0 ) ;
	assign w_sub08_U_r_w = ( (|r_sys_processing_methodID) ? r_sub08_U_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 15'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub24_T_addr = ( (|r_sys_processing_methodID) ? r_sub24_T_addr : 15'sh0 ) ;
	assign w_sub24_T_datain = ( (|r_sys_processing_methodID) ? r_sub24_T_datain : 32'h0 ) ;
	assign w_sub24_T_r_w = ( (|r_sys_processing_methodID) ? r_sub24_T_r_w : 1'h0 ) ;
	assign w_sub24_V_addr = ( (|r_sys_processing_methodID) ? r_sub24_V_addr : 15'sh0 ) ;
	assign w_sub24_V_datain = ( (|r_sys_processing_methodID) ? r_sub24_V_datain : 32'h0 ) ;
	assign w_sub24_V_r_w = ( (|r_sys_processing_methodID) ? r_sub24_V_r_w : 1'h0 ) ;
	assign w_sub24_U_addr = ( (|r_sys_processing_methodID) ? r_sub24_U_addr : 15'sh0 ) ;
	assign w_sub24_U_datain = ( (|r_sys_processing_methodID) ? r_sub24_U_datain : 32'h0 ) ;
	assign w_sub24_U_r_w = ( (|r_sys_processing_methodID) ? r_sub24_U_r_w : 1'h0 ) ;
	assign w_sub24_result_addr = ( (|r_sys_processing_methodID) ? r_sub24_result_addr : 15'sh0 ) ;
	assign w_sub24_result_datain = ( (|r_sys_processing_methodID) ? r_sub24_result_datain : 32'h0 ) ;
	assign w_sub24_result_r_w = ( (|r_sys_processing_methodID) ? r_sub24_result_r_w : 1'h0 ) ;
	assign w_sub25_T_addr = ( (|r_sys_processing_methodID) ? r_sub25_T_addr : 15'sh0 ) ;
	assign w_sub25_T_datain = ( (|r_sys_processing_methodID) ? r_sub25_T_datain : 32'h0 ) ;
	assign w_sub25_T_r_w = ( (|r_sys_processing_methodID) ? r_sub25_T_r_w : 1'h0 ) ;
	assign w_sub25_V_addr = ( (|r_sys_processing_methodID) ? r_sub25_V_addr : 15'sh0 ) ;
	assign w_sub25_V_datain = ( (|r_sys_processing_methodID) ? r_sub25_V_datain : 32'h0 ) ;
	assign w_sub25_V_r_w = ( (|r_sys_processing_methodID) ? r_sub25_V_r_w : 1'h0 ) ;
	assign w_sub25_U_addr = ( (|r_sys_processing_methodID) ? r_sub25_U_addr : 15'sh0 ) ;
	assign w_sub25_U_datain = ( (|r_sys_processing_methodID) ? r_sub25_U_datain : 32'h0 ) ;
	assign w_sub25_U_r_w = ( (|r_sys_processing_methodID) ? r_sub25_U_r_w : 1'h0 ) ;
	assign w_sub25_result_addr = ( (|r_sys_processing_methodID) ? r_sub25_result_addr : 15'sh0 ) ;
	assign w_sub25_result_datain = ( (|r_sys_processing_methodID) ? r_sub25_result_datain : 32'h0 ) ;
	assign w_sub25_result_r_w = ( (|r_sys_processing_methodID) ? r_sub25_result_r_w : 1'h0 ) ;
	assign w_sub22_T_addr = ( (|r_sys_processing_methodID) ? r_sub22_T_addr : 15'sh0 ) ;
	assign w_sub22_T_datain = ( (|r_sys_processing_methodID) ? r_sub22_T_datain : 32'h0 ) ;
	assign w_sub22_T_r_w = ( (|r_sys_processing_methodID) ? r_sub22_T_r_w : 1'h0 ) ;
	assign w_sub22_V_addr = ( (|r_sys_processing_methodID) ? r_sub22_V_addr : 15'sh0 ) ;
	assign w_sub22_V_datain = ( (|r_sys_processing_methodID) ? r_sub22_V_datain : 32'h0 ) ;
	assign w_sub22_V_r_w = ( (|r_sys_processing_methodID) ? r_sub22_V_r_w : 1'h0 ) ;
	assign w_sub22_U_addr = ( (|r_sys_processing_methodID) ? r_sub22_U_addr : 15'sh0 ) ;
	assign w_sub22_U_datain = ( (|r_sys_processing_methodID) ? r_sub22_U_datain : 32'h0 ) ;
	assign w_sub22_U_r_w = ( (|r_sys_processing_methodID) ? r_sub22_U_r_w : 1'h0 ) ;
	assign w_sub22_result_addr = ( (|r_sys_processing_methodID) ? r_sub22_result_addr : 15'sh0 ) ;
	assign w_sub22_result_datain = ( (|r_sys_processing_methodID) ? r_sub22_result_datain : 32'h0 ) ;
	assign w_sub22_result_r_w = ( (|r_sys_processing_methodID) ? r_sub22_result_r_w : 1'h0 ) ;
	assign w_sub23_T_addr = ( (|r_sys_processing_methodID) ? r_sub23_T_addr : 15'sh0 ) ;
	assign w_sub23_T_datain = ( (|r_sys_processing_methodID) ? r_sub23_T_datain : 32'h0 ) ;
	assign w_sub23_T_r_w = ( (|r_sys_processing_methodID) ? r_sub23_T_r_w : 1'h0 ) ;
	assign w_sub23_V_addr = ( (|r_sys_processing_methodID) ? r_sub23_V_addr : 15'sh0 ) ;
	assign w_sub23_V_datain = ( (|r_sys_processing_methodID) ? r_sub23_V_datain : 32'h0 ) ;
	assign w_sub23_V_r_w = ( (|r_sys_processing_methodID) ? r_sub23_V_r_w : 1'h0 ) ;
	assign w_sub23_U_addr = ( (|r_sys_processing_methodID) ? r_sub23_U_addr : 15'sh0 ) ;
	assign w_sub23_U_datain = ( (|r_sys_processing_methodID) ? r_sub23_U_datain : 32'h0 ) ;
	assign w_sub23_U_r_w = ( (|r_sys_processing_methodID) ? r_sub23_U_r_w : 1'h0 ) ;
	assign w_sub23_result_addr = ( (|r_sys_processing_methodID) ? r_sub23_result_addr : 15'sh0 ) ;
	assign w_sub23_result_datain = ( (|r_sys_processing_methodID) ? r_sub23_result_datain : 32'h0 ) ;
	assign w_sub23_result_r_w = ( (|r_sys_processing_methodID) ? r_sub23_result_r_w : 1'h0 ) ;
	assign w_sub03_T_addr = ( (|r_sys_processing_methodID) ? r_sub03_T_addr : 15'sh0 ) ;
	assign w_sub03_T_datain = ( (|r_sys_processing_methodID) ? r_sub03_T_datain : 32'h0 ) ;
	assign w_sub03_T_r_w = ( (|r_sys_processing_methodID) ? r_sub03_T_r_w : 1'h0 ) ;
	assign w_sub03_V_addr = ( (|r_sys_processing_methodID) ? r_sub03_V_addr : 15'sh0 ) ;
	assign w_sub03_V_datain = ( (|r_sys_processing_methodID) ? r_sub03_V_datain : 32'h0 ) ;
	assign w_sub03_V_r_w = ( (|r_sys_processing_methodID) ? r_sub03_V_r_w : 1'h0 ) ;
	assign w_sub03_U_addr = ( (|r_sys_processing_methodID) ? r_sub03_U_addr : 15'sh0 ) ;
	assign w_sub03_U_datain = ( (|r_sys_processing_methodID) ? r_sub03_U_datain : 32'h0 ) ;
	assign w_sub03_U_r_w = ( (|r_sys_processing_methodID) ? r_sub03_U_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 15'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_T_addr = ( (|r_sys_processing_methodID) ? r_sub02_T_addr : 15'sh0 ) ;
	assign w_sub02_T_datain = ( (|r_sys_processing_methodID) ? r_sub02_T_datain : 32'h0 ) ;
	assign w_sub02_T_r_w = ( (|r_sys_processing_methodID) ? r_sub02_T_r_w : 1'h0 ) ;
	assign w_sub02_V_addr = ( (|r_sys_processing_methodID) ? r_sub02_V_addr : 15'sh0 ) ;
	assign w_sub02_V_datain = ( (|r_sys_processing_methodID) ? r_sub02_V_datain : 32'h0 ) ;
	assign w_sub02_V_r_w = ( (|r_sys_processing_methodID) ? r_sub02_V_r_w : 1'h0 ) ;
	assign w_sub02_U_addr = ( (|r_sys_processing_methodID) ? r_sub02_U_addr : 15'sh0 ) ;
	assign w_sub02_U_datain = ( (|r_sys_processing_methodID) ? r_sub02_U_datain : 32'h0 ) ;
	assign w_sub02_U_r_w = ( (|r_sys_processing_methodID) ? r_sub02_U_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 15'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_T_addr = ( (|r_sys_processing_methodID) ? r_sub01_T_addr : 15'sh0 ) ;
	assign w_sub01_T_datain = ( (|r_sys_processing_methodID) ? r_sub01_T_datain : 32'h0 ) ;
	assign w_sub01_T_r_w = ( (|r_sys_processing_methodID) ? r_sub01_T_r_w : 1'h0 ) ;
	assign w_sub01_V_addr = ( (|r_sys_processing_methodID) ? r_sub01_V_addr : 15'sh0 ) ;
	assign w_sub01_V_datain = ( (|r_sys_processing_methodID) ? r_sub01_V_datain : 32'h0 ) ;
	assign w_sub01_V_r_w = ( (|r_sys_processing_methodID) ? r_sub01_V_r_w : 1'h0 ) ;
	assign w_sub01_U_addr = ( (|r_sys_processing_methodID) ? r_sub01_U_addr : 15'sh0 ) ;
	assign w_sub01_U_datain = ( (|r_sys_processing_methodID) ? r_sub01_U_datain : 32'h0 ) ;
	assign w_sub01_U_r_w = ( (|r_sys_processing_methodID) ? r_sub01_U_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 15'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_T_addr = ( (|r_sys_processing_methodID) ? r_sub00_T_addr : 15'sh0 ) ;
	assign w_sub00_T_datain = ( (|r_sys_processing_methodID) ? r_sub00_T_datain : 32'h0 ) ;
	assign w_sub00_T_r_w = ( (|r_sys_processing_methodID) ? r_sub00_T_r_w : 1'h0 ) ;
	assign w_sub00_V_addr = ( (|r_sys_processing_methodID) ? r_sub00_V_addr : 15'sh0 ) ;
	assign w_sub00_V_datain = ( (|r_sys_processing_methodID) ? r_sub00_V_datain : 32'h0 ) ;
	assign w_sub00_V_r_w = ( (|r_sys_processing_methodID) ? r_sub00_V_r_w : 1'h0 ) ;
	assign w_sub00_U_addr = ( (|r_sys_processing_methodID) ? r_sub00_U_addr : 15'sh0 ) ;
	assign w_sub00_U_datain = ( (|r_sys_processing_methodID) ? r_sub00_U_datain : 32'h0 ) ;
	assign w_sub00_U_r_w = ( (|r_sys_processing_methodID) ? r_sub00_U_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 15'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_T_addr = ( (|r_sys_processing_methodID) ? r_sub07_T_addr : 15'sh0 ) ;
	assign w_sub07_T_datain = ( (|r_sys_processing_methodID) ? r_sub07_T_datain : 32'h0 ) ;
	assign w_sub07_T_r_w = ( (|r_sys_processing_methodID) ? r_sub07_T_r_w : 1'h0 ) ;
	assign w_sub07_V_addr = ( (|r_sys_processing_methodID) ? r_sub07_V_addr : 15'sh0 ) ;
	assign w_sub07_V_datain = ( (|r_sys_processing_methodID) ? r_sub07_V_datain : 32'h0 ) ;
	assign w_sub07_V_r_w = ( (|r_sys_processing_methodID) ? r_sub07_V_r_w : 1'h0 ) ;
	assign w_sub07_U_addr = ( (|r_sys_processing_methodID) ? r_sub07_U_addr : 15'sh0 ) ;
	assign w_sub07_U_datain = ( (|r_sys_processing_methodID) ? r_sub07_U_datain : 32'h0 ) ;
	assign w_sub07_U_r_w = ( (|r_sys_processing_methodID) ? r_sub07_U_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 15'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_T_addr = ( (|r_sys_processing_methodID) ? r_sub06_T_addr : 15'sh0 ) ;
	assign w_sub06_T_datain = ( (|r_sys_processing_methodID) ? r_sub06_T_datain : 32'h0 ) ;
	assign w_sub06_T_r_w = ( (|r_sys_processing_methodID) ? r_sub06_T_r_w : 1'h0 ) ;
	assign w_sub06_V_addr = ( (|r_sys_processing_methodID) ? r_sub06_V_addr : 15'sh0 ) ;
	assign w_sub06_V_datain = ( (|r_sys_processing_methodID) ? r_sub06_V_datain : 32'h0 ) ;
	assign w_sub06_V_r_w = ( (|r_sys_processing_methodID) ? r_sub06_V_r_w : 1'h0 ) ;
	assign w_sub06_U_addr = ( (|r_sys_processing_methodID) ? r_sub06_U_addr : 15'sh0 ) ;
	assign w_sub06_U_datain = ( (|r_sys_processing_methodID) ? r_sub06_U_datain : 32'h0 ) ;
	assign w_sub06_U_r_w = ( (|r_sys_processing_methodID) ? r_sub06_U_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 15'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub05_T_addr = ( (|r_sys_processing_methodID) ? r_sub05_T_addr : 15'sh0 ) ;
	assign w_sub05_T_datain = ( (|r_sys_processing_methodID) ? r_sub05_T_datain : 32'h0 ) ;
	assign w_sub05_T_r_w = ( (|r_sys_processing_methodID) ? r_sub05_T_r_w : 1'h0 ) ;
	assign w_sub05_V_addr = ( (|r_sys_processing_methodID) ? r_sub05_V_addr : 15'sh0 ) ;
	assign w_sub05_V_datain = ( (|r_sys_processing_methodID) ? r_sub05_V_datain : 32'h0 ) ;
	assign w_sub05_V_r_w = ( (|r_sys_processing_methodID) ? r_sub05_V_r_w : 1'h0 ) ;
	assign w_sub05_U_addr = ( (|r_sys_processing_methodID) ? r_sub05_U_addr : 15'sh0 ) ;
	assign w_sub05_U_datain = ( (|r_sys_processing_methodID) ? r_sub05_U_datain : 32'h0 ) ;
	assign w_sub05_U_r_w = ( (|r_sys_processing_methodID) ? r_sub05_U_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 15'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_T_addr = ( (|r_sys_processing_methodID) ? r_sub04_T_addr : 15'sh0 ) ;
	assign w_sub04_T_datain = ( (|r_sys_processing_methodID) ? r_sub04_T_datain : 32'h0 ) ;
	assign w_sub04_T_r_w = ( (|r_sys_processing_methodID) ? r_sub04_T_r_w : 1'h0 ) ;
	assign w_sub04_V_addr = ( (|r_sys_processing_methodID) ? r_sub04_V_addr : 15'sh0 ) ;
	assign w_sub04_V_datain = ( (|r_sys_processing_methodID) ? r_sub04_V_datain : 32'h0 ) ;
	assign w_sub04_V_r_w = ( (|r_sys_processing_methodID) ? r_sub04_V_r_w : 1'h0 ) ;
	assign w_sub04_U_addr = ( (|r_sys_processing_methodID) ? r_sub04_U_addr : 15'sh0 ) ;
	assign w_sub04_U_datain = ( (|r_sys_processing_methodID) ? r_sub04_U_datain : 32'h0 ) ;
	assign w_sub04_U_r_w = ( (|r_sys_processing_methodID) ? r_sub04_U_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 15'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_T_addr = ( (|r_sys_processing_methodID) ? r_sub10_T_addr : 15'sh0 ) ;
	assign w_sub10_T_datain = ( (|r_sys_processing_methodID) ? r_sub10_T_datain : 32'h0 ) ;
	assign w_sub10_T_r_w = ( (|r_sys_processing_methodID) ? r_sub10_T_r_w : 1'h0 ) ;
	assign w_sub10_V_addr = ( (|r_sys_processing_methodID) ? r_sub10_V_addr : 15'sh0 ) ;
	assign w_sub10_V_datain = ( (|r_sys_processing_methodID) ? r_sub10_V_datain : 32'h0 ) ;
	assign w_sub10_V_r_w = ( (|r_sys_processing_methodID) ? r_sub10_V_r_w : 1'h0 ) ;
	assign w_sub10_U_addr = ( (|r_sys_processing_methodID) ? r_sub10_U_addr : 15'sh0 ) ;
	assign w_sub10_U_datain = ( (|r_sys_processing_methodID) ? r_sub10_U_datain : 32'h0 ) ;
	assign w_sub10_U_r_w = ( (|r_sys_processing_methodID) ? r_sub10_U_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 15'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sub31_T_addr = ( (|r_sys_processing_methodID) ? r_sub31_T_addr : 15'sh0 ) ;
	assign w_sub31_T_datain = ( (|r_sys_processing_methodID) ? r_sub31_T_datain : 32'h0 ) ;
	assign w_sub31_T_r_w = ( (|r_sys_processing_methodID) ? r_sub31_T_r_w : 1'h0 ) ;
	assign w_sub31_V_addr = ( (|r_sys_processing_methodID) ? r_sub31_V_addr : 15'sh0 ) ;
	assign w_sub31_V_datain = ( (|r_sys_processing_methodID) ? r_sub31_V_datain : 32'h0 ) ;
	assign w_sub31_V_r_w = ( (|r_sys_processing_methodID) ? r_sub31_V_r_w : 1'h0 ) ;
	assign w_sub31_U_addr = ( (|r_sys_processing_methodID) ? r_sub31_U_addr : 15'sh0 ) ;
	assign w_sub31_U_datain = ( (|r_sys_processing_methodID) ? r_sub31_U_datain : 32'h0 ) ;
	assign w_sub31_U_r_w = ( (|r_sys_processing_methodID) ? r_sub31_U_r_w : 1'h0 ) ;
	assign w_sub31_result_addr = ( (|r_sys_processing_methodID) ? r_sub31_result_addr : 15'sh0 ) ;
	assign w_sub31_result_datain = ( (|r_sys_processing_methodID) ? r_sub31_result_datain : 32'h0 ) ;
	assign w_sub31_result_r_w = ( (|r_sys_processing_methodID) ? r_sub31_result_r_w : 1'h0 ) ;
	assign w_sub30_T_addr = ( (|r_sys_processing_methodID) ? r_sub30_T_addr : 15'sh0 ) ;
	assign w_sub30_T_datain = ( (|r_sys_processing_methodID) ? r_sub30_T_datain : 32'h0 ) ;
	assign w_sub30_T_r_w = ( (|r_sys_processing_methodID) ? r_sub30_T_r_w : 1'h0 ) ;
	assign w_sub30_V_addr = ( (|r_sys_processing_methodID) ? r_sub30_V_addr : 15'sh0 ) ;
	assign w_sub30_V_datain = ( (|r_sys_processing_methodID) ? r_sub30_V_datain : 32'h0 ) ;
	assign w_sub30_V_r_w = ( (|r_sys_processing_methodID) ? r_sub30_V_r_w : 1'h0 ) ;
	assign w_sub30_U_addr = ( (|r_sys_processing_methodID) ? r_sub30_U_addr : 15'sh0 ) ;
	assign w_sub30_U_datain = ( (|r_sys_processing_methodID) ? r_sub30_U_datain : 32'h0 ) ;
	assign w_sub30_U_r_w = ( (|r_sys_processing_methodID) ? r_sub30_U_r_w : 1'h0 ) ;
	assign w_sub30_result_addr = ( (|r_sys_processing_methodID) ? r_sub30_result_addr : 15'sh0 ) ;
	assign w_sub30_result_datain = ( (|r_sys_processing_methodID) ? r_sub30_result_datain : 32'h0 ) ;
	assign w_sub30_result_r_w = ( (|r_sys_processing_methodID) ? r_sub30_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000080;
	assign w_sys_tmp3 = 32'sh00000081;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'h3d000000;
	assign w_sys_tmp7 = 32'h3c000000;
	assign w_sys_tmp8 = 32'h3c03126f;
	assign w_sys_tmp9 = 32'h3d03126f;
	assign w_sys_tmp10 = 32'h3f03126f;
	assign w_sys_tmp11 = 32'h4103126f;
	assign w_sys_tmp12 = ( !w_sys_tmp13 );
	assign w_sys_tmp13 = (r_run_my_40 < r_run_k_36);
	assign w_sys_tmp14 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp15 = ( !w_sys_tmp16 );
	assign w_sys_tmp16 = (r_run_mx_39 < r_run_j_37);
	assign w_sys_tmp18 = w_ip_MultFloat_product_0;
	assign w_sys_tmp19 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp20 = (r_run_k_36 - w_sys_intOne);
	assign w_sys_tmp22 = (w_sys_tmp23 + r_run_k_36);
	assign w_sys_tmp23 = (r_run_j_37 * w_sys_tmp24);
	assign w_sys_tmp24 = 32'sh00000081;
	assign w_sys_tmp25 = 32'h0;
	assign w_sys_tmp27 = (w_sys_tmp28 + r_run_k_36);
	assign w_sys_tmp28 = (r_run_copy2_j_55 * w_sys_tmp24);
	assign w_sys_tmp32 = (w_sys_tmp33 + r_run_k_36);
	assign w_sys_tmp33 = (r_run_copy1_j_54 * w_sys_tmp24);
	assign w_sys_tmp36 = 32'h42200000;
	assign w_sys_tmp37 = w_sys_tmp18;
	assign w_sys_tmp38 = 32'h3f800000;
	assign w_sys_tmp41 = (w_sys_tmp42 + r_run_k_36);
	assign w_sys_tmp42 = (r_run_copy0_j_53 * w_sys_tmp24);
	assign w_sys_tmp45 = (r_run_copy0_j_53 + w_sys_intOne);
	assign w_sys_tmp46 = (r_run_copy1_j_54 + w_sys_intOne);
	assign w_sys_tmp47 = (r_run_copy2_j_55 + w_sys_intOne);
	assign w_sys_tmp48 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp128 = r_sys_tmp4_float;
	assign w_sys_tmp226 = ( !w_sys_tmp227 );
	assign w_sys_tmp227 = (w_sys_tmp228 < r_run_k_36);
	assign w_sys_tmp228 = 32'sh00000021;
	assign w_sys_tmp229 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp230 = ( !w_sys_tmp231 );
	assign w_sys_tmp231 = (w_sys_tmp232 < r_run_j_37);
	assign w_sys_tmp232 = 32'sh00000011;
	assign w_sys_tmp235 = (w_sys_tmp236 + r_run_k_36);
	assign w_sys_tmp236 = (r_run_j_37 * w_sys_tmp237);
	assign w_sys_tmp237 = 32'sh00000081;
	assign w_sys_tmp238 = w_fld_U_2_dataout_1;
	assign w_sys_tmp239 = (w_sys_tmp240 + r_run_k_36);
	assign w_sys_tmp240 = (r_run_copy4_j_60 * w_sys_tmp237);
	assign w_sys_tmp243 = (w_sys_tmp244 + r_run_k_36);
	assign w_sys_tmp244 = (r_run_copy3_j_59 * w_sys_tmp237);
	assign w_sys_tmp246 = w_fld_V_3_dataout_1;
	assign w_sys_tmp247 = (w_sys_tmp248 + r_run_k_36);
	assign w_sys_tmp248 = (r_run_copy2_j_58 * w_sys_tmp237);
	assign w_sys_tmp251 = (w_sys_tmp252 + r_run_k_36);
	assign w_sys_tmp252 = (r_run_copy1_j_57 * w_sys_tmp237);
	assign w_sys_tmp254 = w_fld_T_0_dataout_1;
	assign w_sys_tmp255 = (w_sys_tmp256 + r_run_k_36);
	assign w_sys_tmp256 = (r_run_copy0_j_56 * w_sys_tmp237);
	assign w_sys_tmp258 = (r_run_copy0_j_56 + w_sys_intOne);
	assign w_sys_tmp259 = (r_run_copy1_j_57 + w_sys_intOne);
	assign w_sys_tmp260 = (r_run_copy2_j_58 + w_sys_intOne);
	assign w_sys_tmp261 = (r_run_copy3_j_59 + w_sys_intOne);
	assign w_sys_tmp262 = (r_run_copy4_j_60 + w_sys_intOne);
	assign w_sys_tmp263 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp444 = 32'sh00000010;
	assign w_sys_tmp445 = ( !w_sys_tmp446 );
	assign w_sys_tmp446 = (w_sys_tmp447 < r_run_j_37);
	assign w_sys_tmp447 = 32'sh00000021;
	assign w_sys_tmp450 = (w_sys_tmp451 + r_run_k_36);
	assign w_sys_tmp451 = (r_run_j_37 * w_sys_tmp452);
	assign w_sys_tmp452 = 32'sh00000081;
	assign w_sys_tmp453 = w_fld_U_2_dataout_1;
	assign w_sys_tmp454 = (w_sys_tmp455 + r_run_k_36);
	assign w_sys_tmp455 = (r_run_copy4_j_65 * w_sys_tmp452);
	assign w_sys_tmp458 = (w_sys_tmp459 + r_run_k_36);
	assign w_sys_tmp459 = (r_run_copy3_j_64 * w_sys_tmp452);
	assign w_sys_tmp461 = w_fld_V_3_dataout_1;
	assign w_sys_tmp462 = (w_sys_tmp463 + r_run_k_36);
	assign w_sys_tmp463 = (r_run_copy2_j_63 * w_sys_tmp452);
	assign w_sys_tmp466 = (w_sys_tmp467 + r_run_k_36);
	assign w_sys_tmp467 = (r_run_copy1_j_62 * w_sys_tmp452);
	assign w_sys_tmp469 = w_fld_T_0_dataout_1;
	assign w_sys_tmp470 = (w_sys_tmp471 + r_run_k_36);
	assign w_sys_tmp471 = (r_run_copy0_j_61 * w_sys_tmp452);
	assign w_sys_tmp473 = (r_run_copy0_j_61 + w_sys_intOne);
	assign w_sys_tmp474 = (r_run_copy1_j_62 + w_sys_intOne);
	assign w_sys_tmp475 = (r_run_copy2_j_63 + w_sys_intOne);
	assign w_sys_tmp476 = (r_run_copy3_j_64 + w_sys_intOne);
	assign w_sys_tmp477 = (r_run_copy4_j_65 + w_sys_intOne);
	assign w_sys_tmp478 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp659 = 32'sh00000020;
	assign w_sys_tmp660 = ( !w_sys_tmp661 );
	assign w_sys_tmp661 = (w_sys_tmp662 < r_run_j_37);
	assign w_sys_tmp662 = 32'sh00000031;
	assign w_sys_tmp665 = (w_sys_tmp666 + r_run_k_36);
	assign w_sys_tmp666 = (r_run_j_37 * w_sys_tmp667);
	assign w_sys_tmp667 = 32'sh00000081;
	assign w_sys_tmp668 = w_fld_U_2_dataout_1;
	assign w_sys_tmp669 = (w_sys_tmp670 + r_run_k_36);
	assign w_sys_tmp670 = (r_run_copy4_j_70 * w_sys_tmp667);
	assign w_sys_tmp673 = (w_sys_tmp674 + r_run_k_36);
	assign w_sys_tmp674 = (r_run_copy3_j_69 * w_sys_tmp667);
	assign w_sys_tmp676 = w_fld_V_3_dataout_1;
	assign w_sys_tmp677 = (w_sys_tmp678 + r_run_k_36);
	assign w_sys_tmp678 = (r_run_copy2_j_68 * w_sys_tmp667);
	assign w_sys_tmp681 = (w_sys_tmp682 + r_run_k_36);
	assign w_sys_tmp682 = (r_run_copy1_j_67 * w_sys_tmp667);
	assign w_sys_tmp684 = w_fld_T_0_dataout_1;
	assign w_sys_tmp685 = (w_sys_tmp686 + r_run_k_36);
	assign w_sys_tmp686 = (r_run_copy0_j_66 * w_sys_tmp667);
	assign w_sys_tmp688 = (r_run_copy0_j_66 + w_sys_intOne);
	assign w_sys_tmp689 = (r_run_copy1_j_67 + w_sys_intOne);
	assign w_sys_tmp690 = (r_run_copy2_j_68 + w_sys_intOne);
	assign w_sys_tmp691 = (r_run_copy3_j_69 + w_sys_intOne);
	assign w_sys_tmp692 = (r_run_copy4_j_70 + w_sys_intOne);
	assign w_sys_tmp693 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp874 = 32'sh00000030;
	assign w_sys_tmp875 = ( !w_sys_tmp876 );
	assign w_sys_tmp876 = (w_sys_tmp877 < r_run_j_37);
	assign w_sys_tmp877 = 32'sh00000041;
	assign w_sys_tmp880 = (w_sys_tmp881 + r_run_k_36);
	assign w_sys_tmp881 = (r_run_j_37 * w_sys_tmp882);
	assign w_sys_tmp882 = 32'sh00000081;
	assign w_sys_tmp883 = w_fld_U_2_dataout_1;
	assign w_sys_tmp884 = (w_sys_tmp885 + r_run_k_36);
	assign w_sys_tmp885 = (r_run_copy4_j_75 * w_sys_tmp882);
	assign w_sys_tmp888 = (w_sys_tmp889 + r_run_k_36);
	assign w_sys_tmp889 = (r_run_copy3_j_74 * w_sys_tmp882);
	assign w_sys_tmp891 = w_fld_V_3_dataout_1;
	assign w_sys_tmp892 = (w_sys_tmp893 + r_run_k_36);
	assign w_sys_tmp893 = (r_run_copy2_j_73 * w_sys_tmp882);
	assign w_sys_tmp896 = (w_sys_tmp897 + r_run_k_36);
	assign w_sys_tmp897 = (r_run_copy1_j_72 * w_sys_tmp882);
	assign w_sys_tmp899 = w_fld_T_0_dataout_1;
	assign w_sys_tmp900 = (w_sys_tmp901 + r_run_k_36);
	assign w_sys_tmp901 = (r_run_copy0_j_71 * w_sys_tmp882);
	assign w_sys_tmp903 = (r_run_copy0_j_71 + w_sys_intOne);
	assign w_sys_tmp904 = (r_run_copy1_j_72 + w_sys_intOne);
	assign w_sys_tmp905 = (r_run_copy2_j_73 + w_sys_intOne);
	assign w_sys_tmp906 = (r_run_copy3_j_74 + w_sys_intOne);
	assign w_sys_tmp907 = (r_run_copy4_j_75 + w_sys_intOne);
	assign w_sys_tmp908 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp1089 = 32'sh00000040;
	assign w_sys_tmp1090 = ( !w_sys_tmp1091 );
	assign w_sys_tmp1091 = (w_sys_tmp1092 < r_run_j_37);
	assign w_sys_tmp1092 = 32'sh00000051;
	assign w_sys_tmp1095 = (w_sys_tmp1096 + r_run_k_36);
	assign w_sys_tmp1096 = (r_run_j_37 * w_sys_tmp1097);
	assign w_sys_tmp1097 = 32'sh00000081;
	assign w_sys_tmp1098 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1099 = (w_sys_tmp1100 + r_run_k_36);
	assign w_sys_tmp1100 = (r_run_copy4_j_80 * w_sys_tmp1097);
	assign w_sys_tmp1103 = (w_sys_tmp1104 + r_run_k_36);
	assign w_sys_tmp1104 = (r_run_copy3_j_79 * w_sys_tmp1097);
	assign w_sys_tmp1106 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1107 = (w_sys_tmp1108 + r_run_k_36);
	assign w_sys_tmp1108 = (r_run_copy2_j_78 * w_sys_tmp1097);
	assign w_sys_tmp1111 = (w_sys_tmp1112 + r_run_k_36);
	assign w_sys_tmp1112 = (r_run_copy1_j_77 * w_sys_tmp1097);
	assign w_sys_tmp1114 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1115 = (w_sys_tmp1116 + r_run_k_36);
	assign w_sys_tmp1116 = (r_run_copy0_j_76 * w_sys_tmp1097);
	assign w_sys_tmp1118 = (r_run_copy0_j_76 + w_sys_intOne);
	assign w_sys_tmp1119 = (r_run_copy1_j_77 + w_sys_intOne);
	assign w_sys_tmp1120 = (r_run_copy2_j_78 + w_sys_intOne);
	assign w_sys_tmp1121 = (r_run_copy3_j_79 + w_sys_intOne);
	assign w_sys_tmp1122 = (r_run_copy4_j_80 + w_sys_intOne);
	assign w_sys_tmp1123 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp1304 = 32'sh00000050;
	assign w_sys_tmp1305 = ( !w_sys_tmp1306 );
	assign w_sys_tmp1306 = (w_sys_tmp1307 < r_run_j_37);
	assign w_sys_tmp1307 = 32'sh00000061;
	assign w_sys_tmp1310 = (w_sys_tmp1311 + r_run_k_36);
	assign w_sys_tmp1311 = (r_run_j_37 * w_sys_tmp1312);
	assign w_sys_tmp1312 = 32'sh00000081;
	assign w_sys_tmp1313 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1314 = (w_sys_tmp1315 + r_run_k_36);
	assign w_sys_tmp1315 = (r_run_copy4_j_85 * w_sys_tmp1312);
	assign w_sys_tmp1318 = (w_sys_tmp1319 + r_run_k_36);
	assign w_sys_tmp1319 = (r_run_copy3_j_84 * w_sys_tmp1312);
	assign w_sys_tmp1321 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1322 = (w_sys_tmp1323 + r_run_k_36);
	assign w_sys_tmp1323 = (r_run_copy2_j_83 * w_sys_tmp1312);
	assign w_sys_tmp1326 = (w_sys_tmp1327 + r_run_k_36);
	assign w_sys_tmp1327 = (r_run_copy1_j_82 * w_sys_tmp1312);
	assign w_sys_tmp1329 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1330 = (w_sys_tmp1331 + r_run_k_36);
	assign w_sys_tmp1331 = (r_run_copy0_j_81 * w_sys_tmp1312);
	assign w_sys_tmp1333 = (r_run_copy0_j_81 + w_sys_intOne);
	assign w_sys_tmp1334 = (r_run_copy1_j_82 + w_sys_intOne);
	assign w_sys_tmp1335 = (r_run_copy2_j_83 + w_sys_intOne);
	assign w_sys_tmp1336 = (r_run_copy3_j_84 + w_sys_intOne);
	assign w_sys_tmp1337 = (r_run_copy4_j_85 + w_sys_intOne);
	assign w_sys_tmp1338 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp1519 = 32'sh00000060;
	assign w_sys_tmp1520 = ( !w_sys_tmp1521 );
	assign w_sys_tmp1521 = (w_sys_tmp1522 < r_run_j_37);
	assign w_sys_tmp1522 = 32'sh00000071;
	assign w_sys_tmp1525 = (w_sys_tmp1526 + r_run_k_36);
	assign w_sys_tmp1526 = (r_run_j_37 * w_sys_tmp1527);
	assign w_sys_tmp1527 = 32'sh00000081;
	assign w_sys_tmp1528 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1529 = (w_sys_tmp1530 + r_run_k_36);
	assign w_sys_tmp1530 = (r_run_copy4_j_90 * w_sys_tmp1527);
	assign w_sys_tmp1533 = (w_sys_tmp1534 + r_run_k_36);
	assign w_sys_tmp1534 = (r_run_copy3_j_89 * w_sys_tmp1527);
	assign w_sys_tmp1536 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1537 = (w_sys_tmp1538 + r_run_k_36);
	assign w_sys_tmp1538 = (r_run_copy2_j_88 * w_sys_tmp1527);
	assign w_sys_tmp1541 = (w_sys_tmp1542 + r_run_k_36);
	assign w_sys_tmp1542 = (r_run_copy1_j_87 * w_sys_tmp1527);
	assign w_sys_tmp1544 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1545 = (w_sys_tmp1546 + r_run_k_36);
	assign w_sys_tmp1546 = (r_run_copy0_j_86 * w_sys_tmp1527);
	assign w_sys_tmp1548 = (r_run_copy0_j_86 + w_sys_intOne);
	assign w_sys_tmp1549 = (r_run_copy1_j_87 + w_sys_intOne);
	assign w_sys_tmp1550 = (r_run_copy2_j_88 + w_sys_intOne);
	assign w_sys_tmp1551 = (r_run_copy3_j_89 + w_sys_intOne);
	assign w_sys_tmp1552 = (r_run_copy4_j_90 + w_sys_intOne);
	assign w_sys_tmp1553 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp1734 = 32'sh00000070;
	assign w_sys_tmp1735 = ( !w_sys_tmp1736 );
	assign w_sys_tmp1736 = (w_sys_tmp1737 < r_run_j_37);
	assign w_sys_tmp1737 = 32'sh00000081;
	assign w_sys_tmp1740 = (w_sys_tmp1741 + r_run_k_36);
	assign w_sys_tmp1741 = (r_run_j_37 * w_sys_tmp1742);
	assign w_sys_tmp1742 = 32'sh00000081;
	assign w_sys_tmp1743 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1744 = (w_sys_tmp1745 + r_run_k_36);
	assign w_sys_tmp1745 = (r_run_copy4_j_95 * w_sys_tmp1742);
	assign w_sys_tmp1748 = (w_sys_tmp1749 + r_run_k_36);
	assign w_sys_tmp1749 = (r_run_copy3_j_94 * w_sys_tmp1742);
	assign w_sys_tmp1751 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1752 = (w_sys_tmp1753 + r_run_k_36);
	assign w_sys_tmp1753 = (r_run_copy2_j_93 * w_sys_tmp1742);
	assign w_sys_tmp1756 = (w_sys_tmp1757 + r_run_k_36);
	assign w_sys_tmp1757 = (r_run_copy1_j_92 * w_sys_tmp1742);
	assign w_sys_tmp1759 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1760 = (w_sys_tmp1761 + r_run_k_36);
	assign w_sys_tmp1761 = (r_run_copy0_j_91 * w_sys_tmp1742);
	assign w_sys_tmp1763 = (r_run_copy0_j_91 + w_sys_intOne);
	assign w_sys_tmp1764 = (r_run_copy1_j_92 + w_sys_intOne);
	assign w_sys_tmp1765 = (r_run_copy2_j_93 + w_sys_intOne);
	assign w_sys_tmp1766 = (r_run_copy3_j_94 + w_sys_intOne);
	assign w_sys_tmp1767 = (r_run_copy4_j_95 + w_sys_intOne);
	assign w_sys_tmp1768 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp1949 = ( !w_sys_tmp1950 );
	assign w_sys_tmp1950 = (w_sys_tmp1951 < r_run_k_36);
	assign w_sys_tmp1951 = 32'sh00000021;
	assign w_sys_tmp1952 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp1953 = ( !w_sys_tmp1954 );
	assign w_sys_tmp1954 = (w_sys_tmp1955 < r_run_j_37);
	assign w_sys_tmp1955 = 32'sh00000011;
	assign w_sys_tmp1958 = (w_sys_tmp1959 + r_run_k_36);
	assign w_sys_tmp1959 = (r_run_j_37 * w_sys_tmp1960);
	assign w_sys_tmp1960 = 32'sh00000081;
	assign w_sys_tmp1961 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1962 = (w_sys_tmp1963 + r_run_k_36);
	assign w_sys_tmp1963 = (r_run_copy4_j_100 * w_sys_tmp1960);
	assign w_sys_tmp1966 = (w_sys_tmp1967 + r_run_k_36);
	assign w_sys_tmp1967 = (r_run_copy3_j_99 * w_sys_tmp1960);
	assign w_sys_tmp1969 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1970 = (w_sys_tmp1971 + r_run_k_36);
	assign w_sys_tmp1971 = (r_run_copy2_j_98 * w_sys_tmp1960);
	assign w_sys_tmp1974 = (w_sys_tmp1975 + r_run_k_36);
	assign w_sys_tmp1975 = (r_run_copy1_j_97 * w_sys_tmp1960);
	assign w_sys_tmp1977 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1978 = (w_sys_tmp1979 + r_run_k_36);
	assign w_sys_tmp1979 = (r_run_copy0_j_96 * w_sys_tmp1960);
	assign w_sys_tmp1981 = (r_run_copy0_j_96 + w_sys_intOne);
	assign w_sys_tmp1982 = (r_run_copy1_j_97 + w_sys_intOne);
	assign w_sys_tmp1983 = (r_run_copy2_j_98 + w_sys_intOne);
	assign w_sys_tmp1984 = (r_run_copy3_j_99 + w_sys_intOne);
	assign w_sys_tmp1985 = (r_run_copy4_j_100 + w_sys_intOne);
	assign w_sys_tmp1986 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp2167 = 32'sh00000010;
	assign w_sys_tmp2168 = ( !w_sys_tmp2169 );
	assign w_sys_tmp2169 = (w_sys_tmp2170 < r_run_j_37);
	assign w_sys_tmp2170 = 32'sh00000021;
	assign w_sys_tmp2173 = (w_sys_tmp2174 + r_run_k_36);
	assign w_sys_tmp2174 = (r_run_j_37 * w_sys_tmp2175);
	assign w_sys_tmp2175 = 32'sh00000081;
	assign w_sys_tmp2176 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2177 = (w_sys_tmp2178 + r_run_k_36);
	assign w_sys_tmp2178 = (r_run_copy4_j_105 * w_sys_tmp2175);
	assign w_sys_tmp2181 = (w_sys_tmp2182 + r_run_k_36);
	assign w_sys_tmp2182 = (r_run_copy3_j_104 * w_sys_tmp2175);
	assign w_sys_tmp2184 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2185 = (w_sys_tmp2186 + r_run_k_36);
	assign w_sys_tmp2186 = (r_run_copy2_j_103 * w_sys_tmp2175);
	assign w_sys_tmp2189 = (w_sys_tmp2190 + r_run_k_36);
	assign w_sys_tmp2190 = (r_run_copy1_j_102 * w_sys_tmp2175);
	assign w_sys_tmp2192 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2193 = (w_sys_tmp2194 + r_run_k_36);
	assign w_sys_tmp2194 = (r_run_copy0_j_101 * w_sys_tmp2175);
	assign w_sys_tmp2196 = (r_run_copy0_j_101 + w_sys_intOne);
	assign w_sys_tmp2197 = (r_run_copy1_j_102 + w_sys_intOne);
	assign w_sys_tmp2198 = (r_run_copy2_j_103 + w_sys_intOne);
	assign w_sys_tmp2199 = (r_run_copy3_j_104 + w_sys_intOne);
	assign w_sys_tmp2200 = (r_run_copy4_j_105 + w_sys_intOne);
	assign w_sys_tmp2201 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp2382 = 32'sh00000020;
	assign w_sys_tmp2383 = ( !w_sys_tmp2384 );
	assign w_sys_tmp2384 = (w_sys_tmp2385 < r_run_j_37);
	assign w_sys_tmp2385 = 32'sh00000031;
	assign w_sys_tmp2388 = (w_sys_tmp2389 + r_run_k_36);
	assign w_sys_tmp2389 = (r_run_j_37 * w_sys_tmp2390);
	assign w_sys_tmp2390 = 32'sh00000081;
	assign w_sys_tmp2391 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2392 = (w_sys_tmp2393 + r_run_k_36);
	assign w_sys_tmp2393 = (r_run_copy4_j_110 * w_sys_tmp2390);
	assign w_sys_tmp2396 = (w_sys_tmp2397 + r_run_k_36);
	assign w_sys_tmp2397 = (r_run_copy3_j_109 * w_sys_tmp2390);
	assign w_sys_tmp2399 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2400 = (w_sys_tmp2401 + r_run_k_36);
	assign w_sys_tmp2401 = (r_run_copy2_j_108 * w_sys_tmp2390);
	assign w_sys_tmp2404 = (w_sys_tmp2405 + r_run_k_36);
	assign w_sys_tmp2405 = (r_run_copy1_j_107 * w_sys_tmp2390);
	assign w_sys_tmp2407 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2408 = (w_sys_tmp2409 + r_run_k_36);
	assign w_sys_tmp2409 = (r_run_copy0_j_106 * w_sys_tmp2390);
	assign w_sys_tmp2411 = (r_run_copy0_j_106 + w_sys_intOne);
	assign w_sys_tmp2412 = (r_run_copy1_j_107 + w_sys_intOne);
	assign w_sys_tmp2413 = (r_run_copy2_j_108 + w_sys_intOne);
	assign w_sys_tmp2414 = (r_run_copy3_j_109 + w_sys_intOne);
	assign w_sys_tmp2415 = (r_run_copy4_j_110 + w_sys_intOne);
	assign w_sys_tmp2416 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp2597 = 32'sh00000030;
	assign w_sys_tmp2598 = ( !w_sys_tmp2599 );
	assign w_sys_tmp2599 = (w_sys_tmp2600 < r_run_j_37);
	assign w_sys_tmp2600 = 32'sh00000041;
	assign w_sys_tmp2603 = (w_sys_tmp2604 + r_run_k_36);
	assign w_sys_tmp2604 = (r_run_j_37 * w_sys_tmp2605);
	assign w_sys_tmp2605 = 32'sh00000081;
	assign w_sys_tmp2606 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2607 = (w_sys_tmp2608 + r_run_k_36);
	assign w_sys_tmp2608 = (r_run_copy4_j_115 * w_sys_tmp2605);
	assign w_sys_tmp2611 = (w_sys_tmp2612 + r_run_k_36);
	assign w_sys_tmp2612 = (r_run_copy3_j_114 * w_sys_tmp2605);
	assign w_sys_tmp2614 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2615 = (w_sys_tmp2616 + r_run_k_36);
	assign w_sys_tmp2616 = (r_run_copy2_j_113 * w_sys_tmp2605);
	assign w_sys_tmp2619 = (w_sys_tmp2620 + r_run_k_36);
	assign w_sys_tmp2620 = (r_run_copy1_j_112 * w_sys_tmp2605);
	assign w_sys_tmp2622 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2623 = (w_sys_tmp2624 + r_run_k_36);
	assign w_sys_tmp2624 = (r_run_copy0_j_111 * w_sys_tmp2605);
	assign w_sys_tmp2626 = (r_run_copy0_j_111 + w_sys_intOne);
	assign w_sys_tmp2627 = (r_run_copy1_j_112 + w_sys_intOne);
	assign w_sys_tmp2628 = (r_run_copy2_j_113 + w_sys_intOne);
	assign w_sys_tmp2629 = (r_run_copy3_j_114 + w_sys_intOne);
	assign w_sys_tmp2630 = (r_run_copy4_j_115 + w_sys_intOne);
	assign w_sys_tmp2631 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp2812 = 32'sh00000040;
	assign w_sys_tmp2813 = ( !w_sys_tmp2814 );
	assign w_sys_tmp2814 = (w_sys_tmp2815 < r_run_j_37);
	assign w_sys_tmp2815 = 32'sh00000051;
	assign w_sys_tmp2818 = (w_sys_tmp2819 + r_run_k_36);
	assign w_sys_tmp2819 = (r_run_j_37 * w_sys_tmp2820);
	assign w_sys_tmp2820 = 32'sh00000081;
	assign w_sys_tmp2821 = w_fld_U_2_dataout_1;
	assign w_sys_tmp2822 = (w_sys_tmp2823 + r_run_k_36);
	assign w_sys_tmp2823 = (r_run_copy4_j_120 * w_sys_tmp2820);
	assign w_sys_tmp2826 = (w_sys_tmp2827 + r_run_k_36);
	assign w_sys_tmp2827 = (r_run_copy3_j_119 * w_sys_tmp2820);
	assign w_sys_tmp2829 = w_fld_V_3_dataout_1;
	assign w_sys_tmp2830 = (w_sys_tmp2831 + r_run_k_36);
	assign w_sys_tmp2831 = (r_run_copy2_j_118 * w_sys_tmp2820);
	assign w_sys_tmp2834 = (w_sys_tmp2835 + r_run_k_36);
	assign w_sys_tmp2835 = (r_run_copy1_j_117 * w_sys_tmp2820);
	assign w_sys_tmp2837 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2838 = (w_sys_tmp2839 + r_run_k_36);
	assign w_sys_tmp2839 = (r_run_copy0_j_116 * w_sys_tmp2820);
	assign w_sys_tmp2841 = (r_run_copy0_j_116 + w_sys_intOne);
	assign w_sys_tmp2842 = (r_run_copy1_j_117 + w_sys_intOne);
	assign w_sys_tmp2843 = (r_run_copy2_j_118 + w_sys_intOne);
	assign w_sys_tmp2844 = (r_run_copy3_j_119 + w_sys_intOne);
	assign w_sys_tmp2845 = (r_run_copy4_j_120 + w_sys_intOne);
	assign w_sys_tmp2846 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp3027 = 32'sh00000050;
	assign w_sys_tmp3028 = ( !w_sys_tmp3029 );
	assign w_sys_tmp3029 = (w_sys_tmp3030 < r_run_j_37);
	assign w_sys_tmp3030 = 32'sh00000061;
	assign w_sys_tmp3033 = (w_sys_tmp3034 + r_run_k_36);
	assign w_sys_tmp3034 = (r_run_j_37 * w_sys_tmp3035);
	assign w_sys_tmp3035 = 32'sh00000081;
	assign w_sys_tmp3036 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3037 = (w_sys_tmp3038 + r_run_k_36);
	assign w_sys_tmp3038 = (r_run_copy4_j_125 * w_sys_tmp3035);
	assign w_sys_tmp3041 = (w_sys_tmp3042 + r_run_k_36);
	assign w_sys_tmp3042 = (r_run_copy3_j_124 * w_sys_tmp3035);
	assign w_sys_tmp3044 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3045 = (w_sys_tmp3046 + r_run_k_36);
	assign w_sys_tmp3046 = (r_run_copy2_j_123 * w_sys_tmp3035);
	assign w_sys_tmp3049 = (w_sys_tmp3050 + r_run_k_36);
	assign w_sys_tmp3050 = (r_run_copy1_j_122 * w_sys_tmp3035);
	assign w_sys_tmp3052 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3053 = (w_sys_tmp3054 + r_run_k_36);
	assign w_sys_tmp3054 = (r_run_copy0_j_121 * w_sys_tmp3035);
	assign w_sys_tmp3056 = (r_run_copy0_j_121 + w_sys_intOne);
	assign w_sys_tmp3057 = (r_run_copy1_j_122 + w_sys_intOne);
	assign w_sys_tmp3058 = (r_run_copy2_j_123 + w_sys_intOne);
	assign w_sys_tmp3059 = (r_run_copy3_j_124 + w_sys_intOne);
	assign w_sys_tmp3060 = (r_run_copy4_j_125 + w_sys_intOne);
	assign w_sys_tmp3061 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp3242 = 32'sh00000060;
	assign w_sys_tmp3243 = ( !w_sys_tmp3244 );
	assign w_sys_tmp3244 = (w_sys_tmp3245 < r_run_j_37);
	assign w_sys_tmp3245 = 32'sh00000071;
	assign w_sys_tmp3248 = (w_sys_tmp3249 + r_run_k_36);
	assign w_sys_tmp3249 = (r_run_j_37 * w_sys_tmp3250);
	assign w_sys_tmp3250 = 32'sh00000081;
	assign w_sys_tmp3251 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3252 = (w_sys_tmp3253 + r_run_k_36);
	assign w_sys_tmp3253 = (r_run_copy4_j_130 * w_sys_tmp3250);
	assign w_sys_tmp3256 = (w_sys_tmp3257 + r_run_k_36);
	assign w_sys_tmp3257 = (r_run_copy3_j_129 * w_sys_tmp3250);
	assign w_sys_tmp3259 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3260 = (w_sys_tmp3261 + r_run_k_36);
	assign w_sys_tmp3261 = (r_run_copy2_j_128 * w_sys_tmp3250);
	assign w_sys_tmp3264 = (w_sys_tmp3265 + r_run_k_36);
	assign w_sys_tmp3265 = (r_run_copy1_j_127 * w_sys_tmp3250);
	assign w_sys_tmp3267 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3268 = (w_sys_tmp3269 + r_run_k_36);
	assign w_sys_tmp3269 = (r_run_copy0_j_126 * w_sys_tmp3250);
	assign w_sys_tmp3271 = (r_run_copy0_j_126 + w_sys_intOne);
	assign w_sys_tmp3272 = (r_run_copy1_j_127 + w_sys_intOne);
	assign w_sys_tmp3273 = (r_run_copy2_j_128 + w_sys_intOne);
	assign w_sys_tmp3274 = (r_run_copy3_j_129 + w_sys_intOne);
	assign w_sys_tmp3275 = (r_run_copy4_j_130 + w_sys_intOne);
	assign w_sys_tmp3276 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp3457 = 32'sh00000070;
	assign w_sys_tmp3458 = ( !w_sys_tmp3459 );
	assign w_sys_tmp3459 = (w_sys_tmp3460 < r_run_j_37);
	assign w_sys_tmp3460 = 32'sh00000081;
	assign w_sys_tmp3463 = (w_sys_tmp3464 + r_run_k_36);
	assign w_sys_tmp3464 = (r_run_j_37 * w_sys_tmp3465);
	assign w_sys_tmp3465 = 32'sh00000081;
	assign w_sys_tmp3466 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3467 = (w_sys_tmp3468 + r_run_k_36);
	assign w_sys_tmp3468 = (r_run_copy4_j_135 * w_sys_tmp3465);
	assign w_sys_tmp3471 = (w_sys_tmp3472 + r_run_k_36);
	assign w_sys_tmp3472 = (r_run_copy3_j_134 * w_sys_tmp3465);
	assign w_sys_tmp3474 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3475 = (w_sys_tmp3476 + r_run_k_36);
	assign w_sys_tmp3476 = (r_run_copy2_j_133 * w_sys_tmp3465);
	assign w_sys_tmp3479 = (w_sys_tmp3480 + r_run_k_36);
	assign w_sys_tmp3480 = (r_run_copy1_j_132 * w_sys_tmp3465);
	assign w_sys_tmp3482 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3483 = (w_sys_tmp3484 + r_run_k_36);
	assign w_sys_tmp3484 = (r_run_copy0_j_131 * w_sys_tmp3465);
	assign w_sys_tmp3486 = (r_run_copy0_j_131 + w_sys_intOne);
	assign w_sys_tmp3487 = (r_run_copy1_j_132 + w_sys_intOne);
	assign w_sys_tmp3488 = (r_run_copy2_j_133 + w_sys_intOne);
	assign w_sys_tmp3489 = (r_run_copy3_j_134 + w_sys_intOne);
	assign w_sys_tmp3490 = (r_run_copy4_j_135 + w_sys_intOne);
	assign w_sys_tmp3491 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp3672 = ( !w_sys_tmp3673 );
	assign w_sys_tmp3673 = (w_sys_tmp3674 < r_run_k_36);
	assign w_sys_tmp3674 = 32'sh00000021;
	assign w_sys_tmp3675 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp3676 = ( !w_sys_tmp3677 );
	assign w_sys_tmp3677 = (w_sys_tmp3678 < r_run_j_37);
	assign w_sys_tmp3678 = 32'sh00000011;
	assign w_sys_tmp3681 = (w_sys_tmp3682 + r_run_k_36);
	assign w_sys_tmp3682 = (r_run_j_37 * w_sys_tmp3683);
	assign w_sys_tmp3683 = 32'sh00000081;
	assign w_sys_tmp3684 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3685 = (w_sys_tmp3686 + r_run_k_36);
	assign w_sys_tmp3686 = (r_run_copy4_j_140 * w_sys_tmp3683);
	assign w_sys_tmp3689 = (w_sys_tmp3690 + r_run_k_36);
	assign w_sys_tmp3690 = (r_run_copy3_j_139 * w_sys_tmp3683);
	assign w_sys_tmp3692 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3693 = (w_sys_tmp3694 + r_run_k_36);
	assign w_sys_tmp3694 = (r_run_copy2_j_138 * w_sys_tmp3683);
	assign w_sys_tmp3697 = (w_sys_tmp3698 + r_run_k_36);
	assign w_sys_tmp3698 = (r_run_copy1_j_137 * w_sys_tmp3683);
	assign w_sys_tmp3700 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3701 = (w_sys_tmp3702 + r_run_k_36);
	assign w_sys_tmp3702 = (r_run_copy0_j_136 * w_sys_tmp3683);
	assign w_sys_tmp3704 = (r_run_copy0_j_136 + w_sys_intOne);
	assign w_sys_tmp3705 = (r_run_copy1_j_137 + w_sys_intOne);
	assign w_sys_tmp3706 = (r_run_copy2_j_138 + w_sys_intOne);
	assign w_sys_tmp3707 = (r_run_copy3_j_139 + w_sys_intOne);
	assign w_sys_tmp3708 = (r_run_copy4_j_140 + w_sys_intOne);
	assign w_sys_tmp3709 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp3890 = 32'sh00000010;
	assign w_sys_tmp3891 = ( !w_sys_tmp3892 );
	assign w_sys_tmp3892 = (w_sys_tmp3893 < r_run_j_37);
	assign w_sys_tmp3893 = 32'sh00000021;
	assign w_sys_tmp3896 = (w_sys_tmp3897 + r_run_k_36);
	assign w_sys_tmp3897 = (r_run_j_37 * w_sys_tmp3898);
	assign w_sys_tmp3898 = 32'sh00000081;
	assign w_sys_tmp3899 = w_fld_U_2_dataout_1;
	assign w_sys_tmp3900 = (w_sys_tmp3901 + r_run_k_36);
	assign w_sys_tmp3901 = (r_run_copy4_j_145 * w_sys_tmp3898);
	assign w_sys_tmp3904 = (w_sys_tmp3905 + r_run_k_36);
	assign w_sys_tmp3905 = (r_run_copy3_j_144 * w_sys_tmp3898);
	assign w_sys_tmp3907 = w_fld_V_3_dataout_1;
	assign w_sys_tmp3908 = (w_sys_tmp3909 + r_run_k_36);
	assign w_sys_tmp3909 = (r_run_copy2_j_143 * w_sys_tmp3898);
	assign w_sys_tmp3912 = (w_sys_tmp3913 + r_run_k_36);
	assign w_sys_tmp3913 = (r_run_copy1_j_142 * w_sys_tmp3898);
	assign w_sys_tmp3915 = w_fld_T_0_dataout_1;
	assign w_sys_tmp3916 = (w_sys_tmp3917 + r_run_k_36);
	assign w_sys_tmp3917 = (r_run_copy0_j_141 * w_sys_tmp3898);
	assign w_sys_tmp3919 = (r_run_copy0_j_141 + w_sys_intOne);
	assign w_sys_tmp3920 = (r_run_copy1_j_142 + w_sys_intOne);
	assign w_sys_tmp3921 = (r_run_copy2_j_143 + w_sys_intOne);
	assign w_sys_tmp3922 = (r_run_copy3_j_144 + w_sys_intOne);
	assign w_sys_tmp3923 = (r_run_copy4_j_145 + w_sys_intOne);
	assign w_sys_tmp3924 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp4105 = 32'sh00000020;
	assign w_sys_tmp4106 = ( !w_sys_tmp4107 );
	assign w_sys_tmp4107 = (w_sys_tmp4108 < r_run_j_37);
	assign w_sys_tmp4108 = 32'sh00000031;
	assign w_sys_tmp4111 = (w_sys_tmp4112 + r_run_k_36);
	assign w_sys_tmp4112 = (r_run_j_37 * w_sys_tmp4113);
	assign w_sys_tmp4113 = 32'sh00000081;
	assign w_sys_tmp4114 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4115 = (w_sys_tmp4116 + r_run_k_36);
	assign w_sys_tmp4116 = (r_run_copy4_j_150 * w_sys_tmp4113);
	assign w_sys_tmp4119 = (w_sys_tmp4120 + r_run_k_36);
	assign w_sys_tmp4120 = (r_run_copy3_j_149 * w_sys_tmp4113);
	assign w_sys_tmp4122 = w_fld_V_3_dataout_1;
	assign w_sys_tmp4123 = (w_sys_tmp4124 + r_run_k_36);
	assign w_sys_tmp4124 = (r_run_copy2_j_148 * w_sys_tmp4113);
	assign w_sys_tmp4127 = (w_sys_tmp4128 + r_run_k_36);
	assign w_sys_tmp4128 = (r_run_copy1_j_147 * w_sys_tmp4113);
	assign w_sys_tmp4130 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4131 = (w_sys_tmp4132 + r_run_k_36);
	assign w_sys_tmp4132 = (r_run_copy0_j_146 * w_sys_tmp4113);
	assign w_sys_tmp4134 = (r_run_copy0_j_146 + w_sys_intOne);
	assign w_sys_tmp4135 = (r_run_copy1_j_147 + w_sys_intOne);
	assign w_sys_tmp4136 = (r_run_copy2_j_148 + w_sys_intOne);
	assign w_sys_tmp4137 = (r_run_copy3_j_149 + w_sys_intOne);
	assign w_sys_tmp4138 = (r_run_copy4_j_150 + w_sys_intOne);
	assign w_sys_tmp4139 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp4320 = 32'sh00000030;
	assign w_sys_tmp4321 = ( !w_sys_tmp4322 );
	assign w_sys_tmp4322 = (w_sys_tmp4323 < r_run_j_37);
	assign w_sys_tmp4323 = 32'sh00000041;
	assign w_sys_tmp4326 = (w_sys_tmp4327 + r_run_k_36);
	assign w_sys_tmp4327 = (r_run_j_37 * w_sys_tmp4328);
	assign w_sys_tmp4328 = 32'sh00000081;
	assign w_sys_tmp4329 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4330 = (w_sys_tmp4331 + r_run_k_36);
	assign w_sys_tmp4331 = (r_run_copy4_j_155 * w_sys_tmp4328);
	assign w_sys_tmp4334 = (w_sys_tmp4335 + r_run_k_36);
	assign w_sys_tmp4335 = (r_run_copy3_j_154 * w_sys_tmp4328);
	assign w_sys_tmp4337 = w_fld_V_3_dataout_1;
	assign w_sys_tmp4338 = (w_sys_tmp4339 + r_run_k_36);
	assign w_sys_tmp4339 = (r_run_copy2_j_153 * w_sys_tmp4328);
	assign w_sys_tmp4342 = (w_sys_tmp4343 + r_run_k_36);
	assign w_sys_tmp4343 = (r_run_copy1_j_152 * w_sys_tmp4328);
	assign w_sys_tmp4345 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4346 = (w_sys_tmp4347 + r_run_k_36);
	assign w_sys_tmp4347 = (r_run_copy0_j_151 * w_sys_tmp4328);
	assign w_sys_tmp4349 = (r_run_copy0_j_151 + w_sys_intOne);
	assign w_sys_tmp4350 = (r_run_copy1_j_152 + w_sys_intOne);
	assign w_sys_tmp4351 = (r_run_copy2_j_153 + w_sys_intOne);
	assign w_sys_tmp4352 = (r_run_copy3_j_154 + w_sys_intOne);
	assign w_sys_tmp4353 = (r_run_copy4_j_155 + w_sys_intOne);
	assign w_sys_tmp4354 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp4535 = 32'sh00000040;
	assign w_sys_tmp4536 = ( !w_sys_tmp4537 );
	assign w_sys_tmp4537 = (w_sys_tmp4538 < r_run_j_37);
	assign w_sys_tmp4538 = 32'sh00000051;
	assign w_sys_tmp4541 = (w_sys_tmp4542 + r_run_k_36);
	assign w_sys_tmp4542 = (r_run_j_37 * w_sys_tmp4543);
	assign w_sys_tmp4543 = 32'sh00000081;
	assign w_sys_tmp4544 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4545 = (w_sys_tmp4546 + r_run_k_36);
	assign w_sys_tmp4546 = (r_run_copy4_j_160 * w_sys_tmp4543);
	assign w_sys_tmp4549 = (w_sys_tmp4550 + r_run_k_36);
	assign w_sys_tmp4550 = (r_run_copy3_j_159 * w_sys_tmp4543);
	assign w_sys_tmp4552 = w_fld_V_3_dataout_1;
	assign w_sys_tmp4553 = (w_sys_tmp4554 + r_run_k_36);
	assign w_sys_tmp4554 = (r_run_copy2_j_158 * w_sys_tmp4543);
	assign w_sys_tmp4557 = (w_sys_tmp4558 + r_run_k_36);
	assign w_sys_tmp4558 = (r_run_copy1_j_157 * w_sys_tmp4543);
	assign w_sys_tmp4560 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4561 = (w_sys_tmp4562 + r_run_k_36);
	assign w_sys_tmp4562 = (r_run_copy0_j_156 * w_sys_tmp4543);
	assign w_sys_tmp4564 = (r_run_copy0_j_156 + w_sys_intOne);
	assign w_sys_tmp4565 = (r_run_copy1_j_157 + w_sys_intOne);
	assign w_sys_tmp4566 = (r_run_copy2_j_158 + w_sys_intOne);
	assign w_sys_tmp4567 = (r_run_copy3_j_159 + w_sys_intOne);
	assign w_sys_tmp4568 = (r_run_copy4_j_160 + w_sys_intOne);
	assign w_sys_tmp4569 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp4750 = 32'sh00000050;
	assign w_sys_tmp4751 = ( !w_sys_tmp4752 );
	assign w_sys_tmp4752 = (w_sys_tmp4753 < r_run_j_37);
	assign w_sys_tmp4753 = 32'sh00000061;
	assign w_sys_tmp4756 = (w_sys_tmp4757 + r_run_k_36);
	assign w_sys_tmp4757 = (r_run_j_37 * w_sys_tmp4758);
	assign w_sys_tmp4758 = 32'sh00000081;
	assign w_sys_tmp4759 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4760 = (w_sys_tmp4761 + r_run_k_36);
	assign w_sys_tmp4761 = (r_run_copy4_j_165 * w_sys_tmp4758);
	assign w_sys_tmp4764 = (w_sys_tmp4765 + r_run_k_36);
	assign w_sys_tmp4765 = (r_run_copy3_j_164 * w_sys_tmp4758);
	assign w_sys_tmp4767 = w_fld_V_3_dataout_1;
	assign w_sys_tmp4768 = (w_sys_tmp4769 + r_run_k_36);
	assign w_sys_tmp4769 = (r_run_copy2_j_163 * w_sys_tmp4758);
	assign w_sys_tmp4772 = (w_sys_tmp4773 + r_run_k_36);
	assign w_sys_tmp4773 = (r_run_copy1_j_162 * w_sys_tmp4758);
	assign w_sys_tmp4775 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4776 = (w_sys_tmp4777 + r_run_k_36);
	assign w_sys_tmp4777 = (r_run_copy0_j_161 * w_sys_tmp4758);
	assign w_sys_tmp4779 = (r_run_copy0_j_161 + w_sys_intOne);
	assign w_sys_tmp4780 = (r_run_copy1_j_162 + w_sys_intOne);
	assign w_sys_tmp4781 = (r_run_copy2_j_163 + w_sys_intOne);
	assign w_sys_tmp4782 = (r_run_copy3_j_164 + w_sys_intOne);
	assign w_sys_tmp4783 = (r_run_copy4_j_165 + w_sys_intOne);
	assign w_sys_tmp4784 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp4965 = 32'sh00000060;
	assign w_sys_tmp4966 = ( !w_sys_tmp4967 );
	assign w_sys_tmp4967 = (w_sys_tmp4968 < r_run_j_37);
	assign w_sys_tmp4968 = 32'sh00000071;
	assign w_sys_tmp4971 = (w_sys_tmp4972 + r_run_k_36);
	assign w_sys_tmp4972 = (r_run_j_37 * w_sys_tmp4973);
	assign w_sys_tmp4973 = 32'sh00000081;
	assign w_sys_tmp4974 = w_fld_U_2_dataout_1;
	assign w_sys_tmp4975 = (w_sys_tmp4976 + r_run_k_36);
	assign w_sys_tmp4976 = (r_run_copy4_j_170 * w_sys_tmp4973);
	assign w_sys_tmp4979 = (w_sys_tmp4980 + r_run_k_36);
	assign w_sys_tmp4980 = (r_run_copy3_j_169 * w_sys_tmp4973);
	assign w_sys_tmp4982 = w_fld_V_3_dataout_1;
	assign w_sys_tmp4983 = (w_sys_tmp4984 + r_run_k_36);
	assign w_sys_tmp4984 = (r_run_copy2_j_168 * w_sys_tmp4973);
	assign w_sys_tmp4987 = (w_sys_tmp4988 + r_run_k_36);
	assign w_sys_tmp4988 = (r_run_copy1_j_167 * w_sys_tmp4973);
	assign w_sys_tmp4990 = w_fld_T_0_dataout_1;
	assign w_sys_tmp4991 = (w_sys_tmp4992 + r_run_k_36);
	assign w_sys_tmp4992 = (r_run_copy0_j_166 * w_sys_tmp4973);
	assign w_sys_tmp4994 = (r_run_copy0_j_166 + w_sys_intOne);
	assign w_sys_tmp4995 = (r_run_copy1_j_167 + w_sys_intOne);
	assign w_sys_tmp4996 = (r_run_copy2_j_168 + w_sys_intOne);
	assign w_sys_tmp4997 = (r_run_copy3_j_169 + w_sys_intOne);
	assign w_sys_tmp4998 = (r_run_copy4_j_170 + w_sys_intOne);
	assign w_sys_tmp4999 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp5180 = 32'sh00000070;
	assign w_sys_tmp5181 = ( !w_sys_tmp5182 );
	assign w_sys_tmp5182 = (w_sys_tmp5183 < r_run_j_37);
	assign w_sys_tmp5183 = 32'sh00000081;
	assign w_sys_tmp5186 = (w_sys_tmp5187 + r_run_k_36);
	assign w_sys_tmp5187 = (r_run_j_37 * w_sys_tmp5188);
	assign w_sys_tmp5188 = 32'sh00000081;
	assign w_sys_tmp5189 = w_fld_U_2_dataout_1;
	assign w_sys_tmp5190 = (w_sys_tmp5191 + r_run_k_36);
	assign w_sys_tmp5191 = (r_run_copy4_j_175 * w_sys_tmp5188);
	assign w_sys_tmp5194 = (w_sys_tmp5195 + r_run_k_36);
	assign w_sys_tmp5195 = (r_run_copy3_j_174 * w_sys_tmp5188);
	assign w_sys_tmp5197 = w_fld_V_3_dataout_1;
	assign w_sys_tmp5198 = (w_sys_tmp5199 + r_run_k_36);
	assign w_sys_tmp5199 = (r_run_copy2_j_173 * w_sys_tmp5188);
	assign w_sys_tmp5202 = (w_sys_tmp5203 + r_run_k_36);
	assign w_sys_tmp5203 = (r_run_copy1_j_172 * w_sys_tmp5188);
	assign w_sys_tmp5205 = w_fld_T_0_dataout_1;
	assign w_sys_tmp5206 = (w_sys_tmp5207 + r_run_k_36);
	assign w_sys_tmp5207 = (r_run_copy0_j_171 * w_sys_tmp5188);
	assign w_sys_tmp5209 = (r_run_copy0_j_171 + w_sys_intOne);
	assign w_sys_tmp5210 = (r_run_copy1_j_172 + w_sys_intOne);
	assign w_sys_tmp5211 = (r_run_copy2_j_173 + w_sys_intOne);
	assign w_sys_tmp5212 = (r_run_copy3_j_174 + w_sys_intOne);
	assign w_sys_tmp5213 = (r_run_copy4_j_175 + w_sys_intOne);
	assign w_sys_tmp5214 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp5395 = ( !w_sys_tmp5396 );
	assign w_sys_tmp5396 = (w_sys_tmp5397 < r_run_k_36);
	assign w_sys_tmp5397 = 32'sh00000021;
	assign w_sys_tmp5398 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp5399 = ( !w_sys_tmp5400 );
	assign w_sys_tmp5400 = (w_sys_tmp5401 < r_run_j_37);
	assign w_sys_tmp5401 = 32'sh00000011;
	assign w_sys_tmp5404 = (w_sys_tmp5405 + r_run_k_36);
	assign w_sys_tmp5405 = (r_run_j_37 * w_sys_tmp5406);
	assign w_sys_tmp5406 = 32'sh00000081;
	assign w_sys_tmp5407 = w_fld_U_2_dataout_1;
	assign w_sys_tmp5408 = (w_sys_tmp5409 + r_run_k_36);
	assign w_sys_tmp5409 = (r_run_copy4_j_180 * w_sys_tmp5406);
	assign w_sys_tmp5412 = (w_sys_tmp5413 + r_run_k_36);
	assign w_sys_tmp5413 = (r_run_copy3_j_179 * w_sys_tmp5406);
	assign w_sys_tmp5415 = w_fld_V_3_dataout_1;
	assign w_sys_tmp5416 = (w_sys_tmp5417 + r_run_k_36);
	assign w_sys_tmp5417 = (r_run_copy2_j_178 * w_sys_tmp5406);
	assign w_sys_tmp5420 = (w_sys_tmp5421 + r_run_k_36);
	assign w_sys_tmp5421 = (r_run_copy1_j_177 * w_sys_tmp5406);
	assign w_sys_tmp5423 = w_fld_T_0_dataout_1;
	assign w_sys_tmp5424 = (w_sys_tmp5425 + r_run_k_36);
	assign w_sys_tmp5425 = (r_run_copy0_j_176 * w_sys_tmp5406);
	assign w_sys_tmp5427 = (r_run_copy0_j_176 + w_sys_intOne);
	assign w_sys_tmp5428 = (r_run_copy1_j_177 + w_sys_intOne);
	assign w_sys_tmp5429 = (r_run_copy2_j_178 + w_sys_intOne);
	assign w_sys_tmp5430 = (r_run_copy3_j_179 + w_sys_intOne);
	assign w_sys_tmp5431 = (r_run_copy4_j_180 + w_sys_intOne);
	assign w_sys_tmp5432 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp5613 = 32'sh00000010;
	assign w_sys_tmp5614 = ( !w_sys_tmp5615 );
	assign w_sys_tmp5615 = (w_sys_tmp5616 < r_run_j_37);
	assign w_sys_tmp5616 = 32'sh00000021;
	assign w_sys_tmp5619 = (w_sys_tmp5620 + r_run_k_36);
	assign w_sys_tmp5620 = (r_run_j_37 * w_sys_tmp5621);
	assign w_sys_tmp5621 = 32'sh00000081;
	assign w_sys_tmp5622 = w_fld_U_2_dataout_1;
	assign w_sys_tmp5623 = (w_sys_tmp5624 + r_run_k_36);
	assign w_sys_tmp5624 = (r_run_copy4_j_185 * w_sys_tmp5621);
	assign w_sys_tmp5627 = (w_sys_tmp5628 + r_run_k_36);
	assign w_sys_tmp5628 = (r_run_copy3_j_184 * w_sys_tmp5621);
	assign w_sys_tmp5630 = w_fld_V_3_dataout_1;
	assign w_sys_tmp5631 = (w_sys_tmp5632 + r_run_k_36);
	assign w_sys_tmp5632 = (r_run_copy2_j_183 * w_sys_tmp5621);
	assign w_sys_tmp5635 = (w_sys_tmp5636 + r_run_k_36);
	assign w_sys_tmp5636 = (r_run_copy1_j_182 * w_sys_tmp5621);
	assign w_sys_tmp5638 = w_fld_T_0_dataout_1;
	assign w_sys_tmp5639 = (w_sys_tmp5640 + r_run_k_36);
	assign w_sys_tmp5640 = (r_run_copy0_j_181 * w_sys_tmp5621);
	assign w_sys_tmp5642 = (r_run_copy0_j_181 + w_sys_intOne);
	assign w_sys_tmp5643 = (r_run_copy1_j_182 + w_sys_intOne);
	assign w_sys_tmp5644 = (r_run_copy2_j_183 + w_sys_intOne);
	assign w_sys_tmp5645 = (r_run_copy3_j_184 + w_sys_intOne);
	assign w_sys_tmp5646 = (r_run_copy4_j_185 + w_sys_intOne);
	assign w_sys_tmp5647 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp5828 = 32'sh00000020;
	assign w_sys_tmp5829 = ( !w_sys_tmp5830 );
	assign w_sys_tmp5830 = (w_sys_tmp5831 < r_run_j_37);
	assign w_sys_tmp5831 = 32'sh00000031;
	assign w_sys_tmp5834 = (w_sys_tmp5835 + r_run_k_36);
	assign w_sys_tmp5835 = (r_run_j_37 * w_sys_tmp5836);
	assign w_sys_tmp5836 = 32'sh00000081;
	assign w_sys_tmp5837 = w_fld_U_2_dataout_1;
	assign w_sys_tmp5838 = (w_sys_tmp5839 + r_run_k_36);
	assign w_sys_tmp5839 = (r_run_copy4_j_190 * w_sys_tmp5836);
	assign w_sys_tmp5842 = (w_sys_tmp5843 + r_run_k_36);
	assign w_sys_tmp5843 = (r_run_copy3_j_189 * w_sys_tmp5836);
	assign w_sys_tmp5845 = w_fld_V_3_dataout_1;
	assign w_sys_tmp5846 = (w_sys_tmp5847 + r_run_k_36);
	assign w_sys_tmp5847 = (r_run_copy2_j_188 * w_sys_tmp5836);
	assign w_sys_tmp5850 = (w_sys_tmp5851 + r_run_k_36);
	assign w_sys_tmp5851 = (r_run_copy1_j_187 * w_sys_tmp5836);
	assign w_sys_tmp5853 = w_fld_T_0_dataout_1;
	assign w_sys_tmp5854 = (w_sys_tmp5855 + r_run_k_36);
	assign w_sys_tmp5855 = (r_run_copy0_j_186 * w_sys_tmp5836);
	assign w_sys_tmp5857 = (r_run_copy0_j_186 + w_sys_intOne);
	assign w_sys_tmp5858 = (r_run_copy1_j_187 + w_sys_intOne);
	assign w_sys_tmp5859 = (r_run_copy2_j_188 + w_sys_intOne);
	assign w_sys_tmp5860 = (r_run_copy3_j_189 + w_sys_intOne);
	assign w_sys_tmp5861 = (r_run_copy4_j_190 + w_sys_intOne);
	assign w_sys_tmp5862 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp6043 = 32'sh00000030;
	assign w_sys_tmp6044 = ( !w_sys_tmp6045 );
	assign w_sys_tmp6045 = (w_sys_tmp6046 < r_run_j_37);
	assign w_sys_tmp6046 = 32'sh00000041;
	assign w_sys_tmp6049 = (w_sys_tmp6050 + r_run_k_36);
	assign w_sys_tmp6050 = (r_run_j_37 * w_sys_tmp6051);
	assign w_sys_tmp6051 = 32'sh00000081;
	assign w_sys_tmp6052 = w_fld_U_2_dataout_1;
	assign w_sys_tmp6053 = (w_sys_tmp6054 + r_run_k_36);
	assign w_sys_tmp6054 = (r_run_copy4_j_195 * w_sys_tmp6051);
	assign w_sys_tmp6057 = (w_sys_tmp6058 + r_run_k_36);
	assign w_sys_tmp6058 = (r_run_copy3_j_194 * w_sys_tmp6051);
	assign w_sys_tmp6060 = w_fld_V_3_dataout_1;
	assign w_sys_tmp6061 = (w_sys_tmp6062 + r_run_k_36);
	assign w_sys_tmp6062 = (r_run_copy2_j_193 * w_sys_tmp6051);
	assign w_sys_tmp6065 = (w_sys_tmp6066 + r_run_k_36);
	assign w_sys_tmp6066 = (r_run_copy1_j_192 * w_sys_tmp6051);
	assign w_sys_tmp6068 = w_fld_T_0_dataout_1;
	assign w_sys_tmp6069 = (w_sys_tmp6070 + r_run_k_36);
	assign w_sys_tmp6070 = (r_run_copy0_j_191 * w_sys_tmp6051);
	assign w_sys_tmp6072 = (r_run_copy0_j_191 + w_sys_intOne);
	assign w_sys_tmp6073 = (r_run_copy1_j_192 + w_sys_intOne);
	assign w_sys_tmp6074 = (r_run_copy2_j_193 + w_sys_intOne);
	assign w_sys_tmp6075 = (r_run_copy3_j_194 + w_sys_intOne);
	assign w_sys_tmp6076 = (r_run_copy4_j_195 + w_sys_intOne);
	assign w_sys_tmp6077 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp6258 = 32'sh00000040;
	assign w_sys_tmp6259 = ( !w_sys_tmp6260 );
	assign w_sys_tmp6260 = (w_sys_tmp6261 < r_run_j_37);
	assign w_sys_tmp6261 = 32'sh00000051;
	assign w_sys_tmp6264 = (w_sys_tmp6265 + r_run_k_36);
	assign w_sys_tmp6265 = (r_run_j_37 * w_sys_tmp6266);
	assign w_sys_tmp6266 = 32'sh00000081;
	assign w_sys_tmp6267 = w_fld_U_2_dataout_1;
	assign w_sys_tmp6268 = (w_sys_tmp6269 + r_run_k_36);
	assign w_sys_tmp6269 = (r_run_copy4_j_200 * w_sys_tmp6266);
	assign w_sys_tmp6272 = (w_sys_tmp6273 + r_run_k_36);
	assign w_sys_tmp6273 = (r_run_copy3_j_199 * w_sys_tmp6266);
	assign w_sys_tmp6275 = w_fld_V_3_dataout_1;
	assign w_sys_tmp6276 = (w_sys_tmp6277 + r_run_k_36);
	assign w_sys_tmp6277 = (r_run_copy2_j_198 * w_sys_tmp6266);
	assign w_sys_tmp6280 = (w_sys_tmp6281 + r_run_k_36);
	assign w_sys_tmp6281 = (r_run_copy1_j_197 * w_sys_tmp6266);
	assign w_sys_tmp6283 = w_fld_T_0_dataout_1;
	assign w_sys_tmp6284 = (w_sys_tmp6285 + r_run_k_36);
	assign w_sys_tmp6285 = (r_run_copy0_j_196 * w_sys_tmp6266);
	assign w_sys_tmp6287 = (r_run_copy0_j_196 + w_sys_intOne);
	assign w_sys_tmp6288 = (r_run_copy1_j_197 + w_sys_intOne);
	assign w_sys_tmp6289 = (r_run_copy2_j_198 + w_sys_intOne);
	assign w_sys_tmp6290 = (r_run_copy3_j_199 + w_sys_intOne);
	assign w_sys_tmp6291 = (r_run_copy4_j_200 + w_sys_intOne);
	assign w_sys_tmp6292 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp6473 = 32'sh00000050;
	assign w_sys_tmp6474 = ( !w_sys_tmp6475 );
	assign w_sys_tmp6475 = (w_sys_tmp6476 < r_run_j_37);
	assign w_sys_tmp6476 = 32'sh00000061;
	assign w_sys_tmp6479 = (w_sys_tmp6480 + r_run_k_36);
	assign w_sys_tmp6480 = (r_run_j_37 * w_sys_tmp6481);
	assign w_sys_tmp6481 = 32'sh00000081;
	assign w_sys_tmp6482 = w_fld_U_2_dataout_1;
	assign w_sys_tmp6483 = (w_sys_tmp6484 + r_run_k_36);
	assign w_sys_tmp6484 = (r_run_copy4_j_205 * w_sys_tmp6481);
	assign w_sys_tmp6487 = (w_sys_tmp6488 + r_run_k_36);
	assign w_sys_tmp6488 = (r_run_copy3_j_204 * w_sys_tmp6481);
	assign w_sys_tmp6490 = w_fld_V_3_dataout_1;
	assign w_sys_tmp6491 = (w_sys_tmp6492 + r_run_k_36);
	assign w_sys_tmp6492 = (r_run_copy2_j_203 * w_sys_tmp6481);
	assign w_sys_tmp6495 = (w_sys_tmp6496 + r_run_k_36);
	assign w_sys_tmp6496 = (r_run_copy1_j_202 * w_sys_tmp6481);
	assign w_sys_tmp6498 = w_fld_T_0_dataout_1;
	assign w_sys_tmp6499 = (w_sys_tmp6500 + r_run_k_36);
	assign w_sys_tmp6500 = (r_run_copy0_j_201 * w_sys_tmp6481);
	assign w_sys_tmp6502 = (r_run_copy0_j_201 + w_sys_intOne);
	assign w_sys_tmp6503 = (r_run_copy1_j_202 + w_sys_intOne);
	assign w_sys_tmp6504 = (r_run_copy2_j_203 + w_sys_intOne);
	assign w_sys_tmp6505 = (r_run_copy3_j_204 + w_sys_intOne);
	assign w_sys_tmp6506 = (r_run_copy4_j_205 + w_sys_intOne);
	assign w_sys_tmp6507 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp6688 = 32'sh00000060;
	assign w_sys_tmp6689 = ( !w_sys_tmp6690 );
	assign w_sys_tmp6690 = (w_sys_tmp6691 < r_run_j_37);
	assign w_sys_tmp6691 = 32'sh00000071;
	assign w_sys_tmp6694 = (w_sys_tmp6695 + r_run_k_36);
	assign w_sys_tmp6695 = (r_run_j_37 * w_sys_tmp6696);
	assign w_sys_tmp6696 = 32'sh00000081;
	assign w_sys_tmp6697 = w_fld_U_2_dataout_1;
	assign w_sys_tmp6698 = (w_sys_tmp6699 + r_run_k_36);
	assign w_sys_tmp6699 = (r_run_copy4_j_210 * w_sys_tmp6696);
	assign w_sys_tmp6702 = (w_sys_tmp6703 + r_run_k_36);
	assign w_sys_tmp6703 = (r_run_copy3_j_209 * w_sys_tmp6696);
	assign w_sys_tmp6705 = w_fld_V_3_dataout_1;
	assign w_sys_tmp6706 = (w_sys_tmp6707 + r_run_k_36);
	assign w_sys_tmp6707 = (r_run_copy2_j_208 * w_sys_tmp6696);
	assign w_sys_tmp6710 = (w_sys_tmp6711 + r_run_k_36);
	assign w_sys_tmp6711 = (r_run_copy1_j_207 * w_sys_tmp6696);
	assign w_sys_tmp6713 = w_fld_T_0_dataout_1;
	assign w_sys_tmp6714 = (w_sys_tmp6715 + r_run_k_36);
	assign w_sys_tmp6715 = (r_run_copy0_j_206 * w_sys_tmp6696);
	assign w_sys_tmp6717 = (r_run_copy0_j_206 + w_sys_intOne);
	assign w_sys_tmp6718 = (r_run_copy1_j_207 + w_sys_intOne);
	assign w_sys_tmp6719 = (r_run_copy2_j_208 + w_sys_intOne);
	assign w_sys_tmp6720 = (r_run_copy3_j_209 + w_sys_intOne);
	assign w_sys_tmp6721 = (r_run_copy4_j_210 + w_sys_intOne);
	assign w_sys_tmp6722 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp6903 = 32'sh00000070;
	assign w_sys_tmp6904 = ( !w_sys_tmp6905 );
	assign w_sys_tmp6905 = (w_sys_tmp6906 < r_run_j_37);
	assign w_sys_tmp6906 = 32'sh00000081;
	assign w_sys_tmp6909 = (w_sys_tmp6910 + r_run_k_36);
	assign w_sys_tmp6910 = (r_run_j_37 * w_sys_tmp6911);
	assign w_sys_tmp6911 = 32'sh00000081;
	assign w_sys_tmp6912 = w_fld_U_2_dataout_1;
	assign w_sys_tmp6913 = (w_sys_tmp6914 + r_run_k_36);
	assign w_sys_tmp6914 = (r_run_copy4_j_215 * w_sys_tmp6911);
	assign w_sys_tmp6917 = (w_sys_tmp6918 + r_run_k_36);
	assign w_sys_tmp6918 = (r_run_copy3_j_214 * w_sys_tmp6911);
	assign w_sys_tmp6920 = w_fld_V_3_dataout_1;
	assign w_sys_tmp6921 = (w_sys_tmp6922 + r_run_k_36);
	assign w_sys_tmp6922 = (r_run_copy2_j_213 * w_sys_tmp6911);
	assign w_sys_tmp6925 = (w_sys_tmp6926 + r_run_k_36);
	assign w_sys_tmp6926 = (r_run_copy1_j_212 * w_sys_tmp6911);
	assign w_sys_tmp6928 = w_fld_T_0_dataout_1;
	assign w_sys_tmp6929 = (w_sys_tmp6930 + r_run_k_36);
	assign w_sys_tmp6930 = (r_run_copy0_j_211 * w_sys_tmp6911);
	assign w_sys_tmp6932 = (r_run_copy0_j_211 + w_sys_intOne);
	assign w_sys_tmp6933 = (r_run_copy1_j_212 + w_sys_intOne);
	assign w_sys_tmp6934 = (r_run_copy2_j_213 + w_sys_intOne);
	assign w_sys_tmp6935 = (r_run_copy3_j_214 + w_sys_intOne);
	assign w_sys_tmp6936 = (r_run_copy4_j_215 + w_sys_intOne);
	assign w_sys_tmp6937 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp7118 = ( !w_sys_tmp7119 );
	assign w_sys_tmp7119 = (r_run_nlast_51 < r_run_n_38);
	assign w_sys_tmp7120 = (r_run_n_38 + w_sys_intOne);
	assign w_sys_tmp7121 = 32'sh00000002;
	assign w_sys_tmp7122 = ( !w_sys_tmp7123 );
	assign w_sys_tmp7123 = (w_sys_tmp7124 < r_run_k_36);
	assign w_sys_tmp7124 = 32'sh00000020;
	assign w_sys_tmp7127 = (w_sys_tmp7128 + r_run_k_36);
	assign w_sys_tmp7128 = 32'sh00000891;
	assign w_sys_tmp7129 = w_sub01_result_dataout;
	assign w_sys_tmp7130 = (w_sys_tmp7131 + r_run_k_36);
	assign w_sys_tmp7131 = 32'sh00000102;
	assign w_sys_tmp7133 = (w_sys_tmp7134 + r_run_k_36);
	assign w_sys_tmp7134 = 32'sh00000081;
	assign w_sys_tmp7135 = w_sub00_result_dataout;
	assign w_sys_tmp7136 = (w_sys_tmp7137 + r_run_k_36);
	assign w_sys_tmp7137 = 32'sh00000810;
	assign w_sys_tmp7139 = (w_sys_tmp7140 + r_run_k_36);
	assign w_sys_tmp7140 = 32'sh00000912;
	assign w_sys_tmp7157 = w_sub02_result_dataout;
	assign w_sys_tmp7168 = w_sub03_result_dataout;
	assign w_sys_tmp7179 = w_sub04_result_dataout;
	assign w_sys_tmp7190 = w_sub05_result_dataout;
	assign w_sys_tmp7201 = w_sub06_result_dataout;
	assign w_sys_tmp7204 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp7205 = 32'sh00000020;
	assign w_sys_tmp7206 = ( !w_sys_tmp7207 );
	assign w_sys_tmp7207 = (w_sys_tmp7208 < r_run_k_36);
	assign w_sys_tmp7208 = 32'sh00000041;
	assign w_sys_tmp7211 = (w_sys_tmp7212 + r_run_k_36);
	assign w_sys_tmp7212 = 32'sh00000891;
	assign w_sys_tmp7213 = w_sub09_result_dataout;
	assign w_sys_tmp7214 = (w_sys_tmp7215 + r_run_k_36);
	assign w_sys_tmp7215 = 32'sh00000102;
	assign w_sys_tmp7217 = (w_sys_tmp7218 + r_run_k_36);
	assign w_sys_tmp7218 = 32'sh00000081;
	assign w_sys_tmp7219 = w_sub08_result_dataout;
	assign w_sys_tmp7220 = (w_sys_tmp7221 + r_run_k_36);
	assign w_sys_tmp7221 = 32'sh00000810;
	assign w_sys_tmp7223 = (w_sys_tmp7224 + r_run_k_36);
	assign w_sys_tmp7224 = 32'sh00000912;
	assign w_sys_tmp7241 = w_sub10_result_dataout;
	assign w_sys_tmp7252 = w_sub11_result_dataout;
	assign w_sys_tmp7263 = w_sub12_result_dataout;
	assign w_sys_tmp7274 = w_sub13_result_dataout;
	assign w_sys_tmp7285 = w_sub14_result_dataout;
	assign w_sys_tmp7288 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp7289 = 32'sh00000040;
	assign w_sys_tmp7290 = ( !w_sys_tmp7291 );
	assign w_sys_tmp7291 = (w_sys_tmp7292 < r_run_k_36);
	assign w_sys_tmp7292 = 32'sh00000061;
	assign w_sys_tmp7295 = (w_sys_tmp7296 + r_run_k_36);
	assign w_sys_tmp7296 = 32'sh00000891;
	assign w_sys_tmp7297 = w_sub17_result_dataout;
	assign w_sys_tmp7298 = (w_sys_tmp7299 + r_run_k_36);
	assign w_sys_tmp7299 = 32'sh00000102;
	assign w_sys_tmp7301 = (w_sys_tmp7302 + r_run_k_36);
	assign w_sys_tmp7302 = 32'sh00000081;
	assign w_sys_tmp7303 = w_sub16_result_dataout;
	assign w_sys_tmp7304 = (w_sys_tmp7305 + r_run_k_36);
	assign w_sys_tmp7305 = 32'sh00000810;
	assign w_sys_tmp7307 = (w_sys_tmp7308 + r_run_k_36);
	assign w_sys_tmp7308 = 32'sh00000912;
	assign w_sys_tmp7325 = w_sub18_result_dataout;
	assign w_sys_tmp7336 = w_sub19_result_dataout;
	assign w_sys_tmp7347 = w_sub20_result_dataout;
	assign w_sys_tmp7358 = w_sub21_result_dataout;
	assign w_sys_tmp7369 = w_sub22_result_dataout;
	assign w_sys_tmp7372 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp7373 = 32'sh00000060;
	assign w_sys_tmp7374 = ( !w_sys_tmp7375 );
	assign w_sys_tmp7375 = (w_sys_tmp7376 < r_run_k_36);
	assign w_sys_tmp7376 = 32'sh00000081;
	assign w_sys_tmp7379 = (w_sys_tmp7380 + r_run_k_36);
	assign w_sys_tmp7380 = 32'sh00000891;
	assign w_sys_tmp7381 = w_sub25_result_dataout;
	assign w_sys_tmp7382 = (w_sys_tmp7383 + r_run_k_36);
	assign w_sys_tmp7383 = 32'sh00000102;
	assign w_sys_tmp7385 = (w_sys_tmp7386 + r_run_k_36);
	assign w_sys_tmp7386 = 32'sh00000081;
	assign w_sys_tmp7387 = w_sub24_result_dataout;
	assign w_sys_tmp7388 = (w_sys_tmp7389 + r_run_k_36);
	assign w_sys_tmp7389 = 32'sh00000810;
	assign w_sys_tmp7391 = (w_sys_tmp7392 + r_run_k_36);
	assign w_sys_tmp7392 = 32'sh00000912;
	assign w_sys_tmp7409 = w_sub26_result_dataout;
	assign w_sys_tmp7420 = w_sub27_result_dataout;
	assign w_sys_tmp7431 = w_sub28_result_dataout;
	assign w_sys_tmp7442 = w_sub29_result_dataout;
	assign w_sys_tmp7453 = w_sub30_result_dataout;
	assign w_sys_tmp7456 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp7457 = ( !w_sys_tmp7458 );
	assign w_sys_tmp7458 = (w_sys_tmp7459 < r_run_j_37);
	assign w_sys_tmp7459 = 32'sh00000011;
	assign w_sys_tmp7462 = (w_sys_tmp7463 + w_sys_tmp7465);
	assign w_sys_tmp7463 = (r_run_j_37 * w_sys_tmp7464);
	assign w_sys_tmp7464 = 32'sh00000081;
	assign w_sys_tmp7465 = 32'sh00000021;
	assign w_sys_tmp7466 = w_sub08_result_dataout;
	assign w_sys_tmp7467 = (w_sys_tmp7468 + w_sys_tmp7465);
	assign w_sys_tmp7468 = (r_run_copy10_j_226 * w_sys_tmp7464);
	assign w_sys_tmp7472 = (w_sys_tmp7473 + w_sys_tmp7475);
	assign w_sys_tmp7473 = (r_run_copy9_j_225 * w_sys_tmp7464);
	assign w_sys_tmp7475 = 32'sh00000020;
	assign w_sys_tmp7476 = w_sub00_result_dataout;
	assign w_sys_tmp7477 = (w_sys_tmp7478 + w_sys_tmp7475);
	assign w_sys_tmp7478 = (r_run_copy8_j_224 * w_sys_tmp7464);
	assign w_sys_tmp7482 = (w_sys_tmp7483 + w_sys_tmp7485);
	assign w_sys_tmp7483 = (r_run_copy7_j_223 * w_sys_tmp7464);
	assign w_sys_tmp7485 = 32'sh00000041;
	assign w_sys_tmp7486 = (w_sys_tmp7487 + w_sys_tmp7485);
	assign w_sys_tmp7487 = (r_run_copy6_j_222 * w_sys_tmp7464);
	assign w_sys_tmp7491 = (w_sys_tmp7492 + w_sys_tmp7494);
	assign w_sys_tmp7492 = (r_run_copy5_j_221 * w_sys_tmp7464);
	assign w_sys_tmp7494 = 32'sh00000040;
	assign w_sys_tmp7496 = (w_sys_tmp7497 + w_sys_tmp7494);
	assign w_sys_tmp7497 = (r_run_copy4_j_220 * w_sys_tmp7464);
	assign w_sys_tmp7501 = (w_sys_tmp7502 + w_sys_tmp7504);
	assign w_sys_tmp7502 = (r_run_copy3_j_219 * w_sys_tmp7464);
	assign w_sys_tmp7504 = 32'sh00000061;
	assign w_sys_tmp7505 = (w_sys_tmp7506 + w_sys_tmp7504);
	assign w_sys_tmp7506 = (r_run_copy2_j_218 * w_sys_tmp7464);
	assign w_sys_tmp7510 = (w_sys_tmp7511 + w_sys_tmp7513);
	assign w_sys_tmp7511 = (r_run_copy1_j_217 * w_sys_tmp7464);
	assign w_sys_tmp7513 = 32'sh00000060;
	assign w_sys_tmp7514 = w_sub16_result_dataout;
	assign w_sys_tmp7515 = (w_sys_tmp7516 + w_sys_tmp7513);
	assign w_sys_tmp7516 = (r_run_copy0_j_216 * w_sys_tmp7464);
	assign w_sys_tmp7519 = (r_run_copy0_j_216 + w_sys_intOne);
	assign w_sys_tmp7520 = (r_run_copy1_j_217 + w_sys_intOne);
	assign w_sys_tmp7521 = (r_run_copy2_j_218 + w_sys_intOne);
	assign w_sys_tmp7522 = (r_run_copy3_j_219 + w_sys_intOne);
	assign w_sys_tmp7523 = (r_run_copy4_j_220 + w_sys_intOne);
	assign w_sys_tmp7524 = (r_run_copy5_j_221 + w_sys_intOne);
	assign w_sys_tmp7525 = (r_run_copy6_j_222 + w_sys_intOne);
	assign w_sys_tmp7526 = (r_run_copy7_j_223 + w_sys_intOne);
	assign w_sys_tmp7527 = (r_run_copy8_j_224 + w_sys_intOne);
	assign w_sys_tmp7528 = (r_run_copy9_j_225 + w_sys_intOne);
	assign w_sys_tmp7529 = (r_run_copy10_j_226 + w_sys_intOne);
	assign w_sys_tmp7530 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp7957 = 32'sh00000010;
	assign w_sys_tmp7958 = ( !w_sys_tmp7959 );
	assign w_sys_tmp7959 = (w_sys_tmp7960 < r_run_j_37);
	assign w_sys_tmp7960 = 32'sh00000021;
	assign w_sys_tmp7963 = (w_sys_tmp7964 + w_sys_tmp7966);
	assign w_sys_tmp7964 = (r_run_j_37 * w_sys_tmp7965);
	assign w_sys_tmp7965 = 32'sh00000081;
	assign w_sys_tmp7966 = 32'sh00000021;
	assign w_sys_tmp7967 = w_sub09_result_dataout;
	assign w_sys_tmp7968 = (w_sys_tmp7969 + w_sys_tmp7966);
	assign w_sys_tmp7969 = (r_run_copy10_j_237 * w_sys_tmp7965);
	assign w_sys_tmp7973 = (w_sys_tmp7974 + w_sys_tmp7976);
	assign w_sys_tmp7974 = (r_run_copy9_j_236 * w_sys_tmp7965);
	assign w_sys_tmp7976 = 32'sh00000020;
	assign w_sys_tmp7977 = w_sub01_result_dataout;
	assign w_sys_tmp7978 = (w_sys_tmp7979 + w_sys_tmp7976);
	assign w_sys_tmp7979 = (r_run_copy8_j_235 * w_sys_tmp7965);
	assign w_sys_tmp7983 = (w_sys_tmp7984 + w_sys_tmp7986);
	assign w_sys_tmp7984 = (r_run_copy7_j_234 * w_sys_tmp7965);
	assign w_sys_tmp7986 = 32'sh00000041;
	assign w_sys_tmp7987 = (w_sys_tmp7988 + w_sys_tmp7986);
	assign w_sys_tmp7988 = (r_run_copy6_j_233 * w_sys_tmp7965);
	assign w_sys_tmp7992 = (w_sys_tmp7993 + w_sys_tmp7995);
	assign w_sys_tmp7993 = (r_run_copy5_j_232 * w_sys_tmp7965);
	assign w_sys_tmp7995 = 32'sh00000040;
	assign w_sys_tmp7997 = (w_sys_tmp7998 + w_sys_tmp7995);
	assign w_sys_tmp7998 = (r_run_copy4_j_231 * w_sys_tmp7965);
	assign w_sys_tmp8002 = (w_sys_tmp8003 + w_sys_tmp8005);
	assign w_sys_tmp8003 = (r_run_copy3_j_230 * w_sys_tmp7965);
	assign w_sys_tmp8005 = 32'sh00000061;
	assign w_sys_tmp8006 = (w_sys_tmp8007 + w_sys_tmp8005);
	assign w_sys_tmp8007 = (r_run_copy2_j_229 * w_sys_tmp7965);
	assign w_sys_tmp8011 = (w_sys_tmp8012 + w_sys_tmp8014);
	assign w_sys_tmp8012 = (r_run_copy1_j_228 * w_sys_tmp7965);
	assign w_sys_tmp8014 = 32'sh00000060;
	assign w_sys_tmp8015 = w_sub17_result_dataout;
	assign w_sys_tmp8016 = (w_sys_tmp8017 + w_sys_tmp8014);
	assign w_sys_tmp8017 = (r_run_copy0_j_227 * w_sys_tmp7965);
	assign w_sys_tmp8020 = (r_run_copy0_j_227 + w_sys_intOne);
	assign w_sys_tmp8021 = (r_run_copy1_j_228 + w_sys_intOne);
	assign w_sys_tmp8022 = (r_run_copy2_j_229 + w_sys_intOne);
	assign w_sys_tmp8023 = (r_run_copy3_j_230 + w_sys_intOne);
	assign w_sys_tmp8024 = (r_run_copy4_j_231 + w_sys_intOne);
	assign w_sys_tmp8025 = (r_run_copy5_j_232 + w_sys_intOne);
	assign w_sys_tmp8026 = (r_run_copy6_j_233 + w_sys_intOne);
	assign w_sys_tmp8027 = (r_run_copy7_j_234 + w_sys_intOne);
	assign w_sys_tmp8028 = (r_run_copy8_j_235 + w_sys_intOne);
	assign w_sys_tmp8029 = (r_run_copy9_j_236 + w_sys_intOne);
	assign w_sys_tmp8030 = (r_run_copy10_j_237 + w_sys_intOne);
	assign w_sys_tmp8031 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp8458 = 32'sh00000020;
	assign w_sys_tmp8459 = ( !w_sys_tmp8460 );
	assign w_sys_tmp8460 = (w_sys_tmp8461 < r_run_j_37);
	assign w_sys_tmp8461 = 32'sh00000031;
	assign w_sys_tmp8464 = (w_sys_tmp8465 + w_sys_tmp8467);
	assign w_sys_tmp8465 = (r_run_j_37 * w_sys_tmp8466);
	assign w_sys_tmp8466 = 32'sh00000081;
	assign w_sys_tmp8467 = 32'sh00000021;
	assign w_sys_tmp8468 = w_sub10_result_dataout;
	assign w_sys_tmp8469 = (w_sys_tmp8470 + w_sys_tmp8467);
	assign w_sys_tmp8470 = (r_run_copy10_j_248 * w_sys_tmp8466);
	assign w_sys_tmp8474 = (w_sys_tmp8475 + w_sys_tmp8477);
	assign w_sys_tmp8475 = (r_run_copy9_j_247 * w_sys_tmp8466);
	assign w_sys_tmp8477 = 32'sh00000020;
	assign w_sys_tmp8478 = w_sub02_result_dataout;
	assign w_sys_tmp8479 = (w_sys_tmp8480 + w_sys_tmp8477);
	assign w_sys_tmp8480 = (r_run_copy8_j_246 * w_sys_tmp8466);
	assign w_sys_tmp8484 = (w_sys_tmp8485 + w_sys_tmp8487);
	assign w_sys_tmp8485 = (r_run_copy7_j_245 * w_sys_tmp8466);
	assign w_sys_tmp8487 = 32'sh00000041;
	assign w_sys_tmp8488 = (w_sys_tmp8489 + w_sys_tmp8487);
	assign w_sys_tmp8489 = (r_run_copy6_j_244 * w_sys_tmp8466);
	assign w_sys_tmp8493 = (w_sys_tmp8494 + w_sys_tmp8496);
	assign w_sys_tmp8494 = (r_run_copy5_j_243 * w_sys_tmp8466);
	assign w_sys_tmp8496 = 32'sh00000040;
	assign w_sys_tmp8498 = (w_sys_tmp8499 + w_sys_tmp8496);
	assign w_sys_tmp8499 = (r_run_copy4_j_242 * w_sys_tmp8466);
	assign w_sys_tmp8503 = (w_sys_tmp8504 + w_sys_tmp8506);
	assign w_sys_tmp8504 = (r_run_copy3_j_241 * w_sys_tmp8466);
	assign w_sys_tmp8506 = 32'sh00000061;
	assign w_sys_tmp8507 = (w_sys_tmp8508 + w_sys_tmp8506);
	assign w_sys_tmp8508 = (r_run_copy2_j_240 * w_sys_tmp8466);
	assign w_sys_tmp8512 = (w_sys_tmp8513 + w_sys_tmp8515);
	assign w_sys_tmp8513 = (r_run_copy1_j_239 * w_sys_tmp8466);
	assign w_sys_tmp8515 = 32'sh00000060;
	assign w_sys_tmp8516 = w_sub18_result_dataout;
	assign w_sys_tmp8517 = (w_sys_tmp8518 + w_sys_tmp8515);
	assign w_sys_tmp8518 = (r_run_copy0_j_238 * w_sys_tmp8466);
	assign w_sys_tmp8521 = (r_run_copy0_j_238 + w_sys_intOne);
	assign w_sys_tmp8522 = (r_run_copy1_j_239 + w_sys_intOne);
	assign w_sys_tmp8523 = (r_run_copy2_j_240 + w_sys_intOne);
	assign w_sys_tmp8524 = (r_run_copy3_j_241 + w_sys_intOne);
	assign w_sys_tmp8525 = (r_run_copy4_j_242 + w_sys_intOne);
	assign w_sys_tmp8526 = (r_run_copy5_j_243 + w_sys_intOne);
	assign w_sys_tmp8527 = (r_run_copy6_j_244 + w_sys_intOne);
	assign w_sys_tmp8528 = (r_run_copy7_j_245 + w_sys_intOne);
	assign w_sys_tmp8529 = (r_run_copy8_j_246 + w_sys_intOne);
	assign w_sys_tmp8530 = (r_run_copy9_j_247 + w_sys_intOne);
	assign w_sys_tmp8531 = (r_run_copy10_j_248 + w_sys_intOne);
	assign w_sys_tmp8532 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp8959 = 32'sh00000030;
	assign w_sys_tmp8960 = ( !w_sys_tmp8961 );
	assign w_sys_tmp8961 = (w_sys_tmp8962 < r_run_j_37);
	assign w_sys_tmp8962 = 32'sh00000041;
	assign w_sys_tmp8965 = (w_sys_tmp8966 + w_sys_tmp8968);
	assign w_sys_tmp8966 = (r_run_j_37 * w_sys_tmp8967);
	assign w_sys_tmp8967 = 32'sh00000081;
	assign w_sys_tmp8968 = 32'sh00000021;
	assign w_sys_tmp8969 = w_sub11_result_dataout;
	assign w_sys_tmp8970 = (w_sys_tmp8971 + w_sys_tmp8968);
	assign w_sys_tmp8971 = (r_run_copy10_j_259 * w_sys_tmp8967);
	assign w_sys_tmp8975 = (w_sys_tmp8976 + w_sys_tmp8978);
	assign w_sys_tmp8976 = (r_run_copy9_j_258 * w_sys_tmp8967);
	assign w_sys_tmp8978 = 32'sh00000020;
	assign w_sys_tmp8979 = w_sub03_result_dataout;
	assign w_sys_tmp8980 = (w_sys_tmp8981 + w_sys_tmp8978);
	assign w_sys_tmp8981 = (r_run_copy8_j_257 * w_sys_tmp8967);
	assign w_sys_tmp8985 = (w_sys_tmp8986 + w_sys_tmp8988);
	assign w_sys_tmp8986 = (r_run_copy7_j_256 * w_sys_tmp8967);
	assign w_sys_tmp8988 = 32'sh00000041;
	assign w_sys_tmp8989 = (w_sys_tmp8990 + w_sys_tmp8988);
	assign w_sys_tmp8990 = (r_run_copy6_j_255 * w_sys_tmp8967);
	assign w_sys_tmp8994 = (w_sys_tmp8995 + w_sys_tmp8997);
	assign w_sys_tmp8995 = (r_run_copy5_j_254 * w_sys_tmp8967);
	assign w_sys_tmp8997 = 32'sh00000040;
	assign w_sys_tmp8999 = (w_sys_tmp9000 + w_sys_tmp8997);
	assign w_sys_tmp9000 = (r_run_copy4_j_253 * w_sys_tmp8967);
	assign w_sys_tmp9004 = (w_sys_tmp9005 + w_sys_tmp9007);
	assign w_sys_tmp9005 = (r_run_copy3_j_252 * w_sys_tmp8967);
	assign w_sys_tmp9007 = 32'sh00000061;
	assign w_sys_tmp9008 = (w_sys_tmp9009 + w_sys_tmp9007);
	assign w_sys_tmp9009 = (r_run_copy2_j_251 * w_sys_tmp8967);
	assign w_sys_tmp9013 = (w_sys_tmp9014 + w_sys_tmp9016);
	assign w_sys_tmp9014 = (r_run_copy1_j_250 * w_sys_tmp8967);
	assign w_sys_tmp9016 = 32'sh00000060;
	assign w_sys_tmp9017 = w_sub19_result_dataout;
	assign w_sys_tmp9018 = (w_sys_tmp9019 + w_sys_tmp9016);
	assign w_sys_tmp9019 = (r_run_copy0_j_249 * w_sys_tmp8967);
	assign w_sys_tmp9022 = (r_run_copy0_j_249 + w_sys_intOne);
	assign w_sys_tmp9023 = (r_run_copy1_j_250 + w_sys_intOne);
	assign w_sys_tmp9024 = (r_run_copy2_j_251 + w_sys_intOne);
	assign w_sys_tmp9025 = (r_run_copy3_j_252 + w_sys_intOne);
	assign w_sys_tmp9026 = (r_run_copy4_j_253 + w_sys_intOne);
	assign w_sys_tmp9027 = (r_run_copy5_j_254 + w_sys_intOne);
	assign w_sys_tmp9028 = (r_run_copy6_j_255 + w_sys_intOne);
	assign w_sys_tmp9029 = (r_run_copy7_j_256 + w_sys_intOne);
	assign w_sys_tmp9030 = (r_run_copy8_j_257 + w_sys_intOne);
	assign w_sys_tmp9031 = (r_run_copy9_j_258 + w_sys_intOne);
	assign w_sys_tmp9032 = (r_run_copy10_j_259 + w_sys_intOne);
	assign w_sys_tmp9033 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp9460 = 32'sh00000040;
	assign w_sys_tmp9461 = ( !w_sys_tmp9462 );
	assign w_sys_tmp9462 = (w_sys_tmp9463 < r_run_j_37);
	assign w_sys_tmp9463 = 32'sh00000051;
	assign w_sys_tmp9466 = (w_sys_tmp9467 + w_sys_tmp9469);
	assign w_sys_tmp9467 = (r_run_j_37 * w_sys_tmp9468);
	assign w_sys_tmp9468 = 32'sh00000081;
	assign w_sys_tmp9469 = 32'sh00000021;
	assign w_sys_tmp9470 = w_sub12_result_dataout;
	assign w_sys_tmp9471 = (w_sys_tmp9472 + w_sys_tmp9469);
	assign w_sys_tmp9472 = (r_run_copy10_j_270 * w_sys_tmp9468);
	assign w_sys_tmp9476 = (w_sys_tmp9477 + w_sys_tmp9479);
	assign w_sys_tmp9477 = (r_run_copy9_j_269 * w_sys_tmp9468);
	assign w_sys_tmp9479 = 32'sh00000020;
	assign w_sys_tmp9480 = w_sub04_result_dataout;
	assign w_sys_tmp9481 = (w_sys_tmp9482 + w_sys_tmp9479);
	assign w_sys_tmp9482 = (r_run_copy8_j_268 * w_sys_tmp9468);
	assign w_sys_tmp9486 = (w_sys_tmp9487 + w_sys_tmp9489);
	assign w_sys_tmp9487 = (r_run_copy7_j_267 * w_sys_tmp9468);
	assign w_sys_tmp9489 = 32'sh00000041;
	assign w_sys_tmp9490 = (w_sys_tmp9491 + w_sys_tmp9489);
	assign w_sys_tmp9491 = (r_run_copy6_j_266 * w_sys_tmp9468);
	assign w_sys_tmp9495 = (w_sys_tmp9496 + w_sys_tmp9498);
	assign w_sys_tmp9496 = (r_run_copy5_j_265 * w_sys_tmp9468);
	assign w_sys_tmp9498 = 32'sh00000040;
	assign w_sys_tmp9500 = (w_sys_tmp9501 + w_sys_tmp9498);
	assign w_sys_tmp9501 = (r_run_copy4_j_264 * w_sys_tmp9468);
	assign w_sys_tmp9505 = (w_sys_tmp9506 + w_sys_tmp9508);
	assign w_sys_tmp9506 = (r_run_copy3_j_263 * w_sys_tmp9468);
	assign w_sys_tmp9508 = 32'sh00000061;
	assign w_sys_tmp9509 = (w_sys_tmp9510 + w_sys_tmp9508);
	assign w_sys_tmp9510 = (r_run_copy2_j_262 * w_sys_tmp9468);
	assign w_sys_tmp9514 = (w_sys_tmp9515 + w_sys_tmp9517);
	assign w_sys_tmp9515 = (r_run_copy1_j_261 * w_sys_tmp9468);
	assign w_sys_tmp9517 = 32'sh00000060;
	assign w_sys_tmp9518 = w_sub20_result_dataout;
	assign w_sys_tmp9519 = (w_sys_tmp9520 + w_sys_tmp9517);
	assign w_sys_tmp9520 = (r_run_copy0_j_260 * w_sys_tmp9468);
	assign w_sys_tmp9523 = (r_run_copy0_j_260 + w_sys_intOne);
	assign w_sys_tmp9524 = (r_run_copy1_j_261 + w_sys_intOne);
	assign w_sys_tmp9525 = (r_run_copy2_j_262 + w_sys_intOne);
	assign w_sys_tmp9526 = (r_run_copy3_j_263 + w_sys_intOne);
	assign w_sys_tmp9527 = (r_run_copy4_j_264 + w_sys_intOne);
	assign w_sys_tmp9528 = (r_run_copy5_j_265 + w_sys_intOne);
	assign w_sys_tmp9529 = (r_run_copy6_j_266 + w_sys_intOne);
	assign w_sys_tmp9530 = (r_run_copy7_j_267 + w_sys_intOne);
	assign w_sys_tmp9531 = (r_run_copy8_j_268 + w_sys_intOne);
	assign w_sys_tmp9532 = (r_run_copy9_j_269 + w_sys_intOne);
	assign w_sys_tmp9533 = (r_run_copy10_j_270 + w_sys_intOne);
	assign w_sys_tmp9534 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp9961 = 32'sh00000050;
	assign w_sys_tmp9962 = ( !w_sys_tmp9963 );
	assign w_sys_tmp9963 = (w_sys_tmp9964 < r_run_j_37);
	assign w_sys_tmp9964 = 32'sh00000061;
	assign w_sys_tmp9967 = (w_sys_tmp9968 + w_sys_tmp9970);
	assign w_sys_tmp9968 = (r_run_j_37 * w_sys_tmp9969);
	assign w_sys_tmp9969 = 32'sh00000081;
	assign w_sys_tmp9970 = 32'sh00000021;
	assign w_sys_tmp9971 = w_sub13_result_dataout;
	assign w_sys_tmp9972 = (w_sys_tmp9973 + w_sys_tmp9970);
	assign w_sys_tmp9973 = (r_run_copy10_j_281 * w_sys_tmp9969);
	assign w_sys_tmp9977 = (w_sys_tmp9978 + w_sys_tmp9980);
	assign w_sys_tmp9978 = (r_run_copy9_j_280 * w_sys_tmp9969);
	assign w_sys_tmp9980 = 32'sh00000020;
	assign w_sys_tmp9981 = w_sub05_result_dataout;
	assign w_sys_tmp9982 = (w_sys_tmp9983 + w_sys_tmp9980);
	assign w_sys_tmp9983 = (r_run_copy8_j_279 * w_sys_tmp9969);
	assign w_sys_tmp9987 = (w_sys_tmp9988 + w_sys_tmp9990);
	assign w_sys_tmp9988 = (r_run_copy7_j_278 * w_sys_tmp9969);
	assign w_sys_tmp9990 = 32'sh00000041;
	assign w_sys_tmp9991 = (w_sys_tmp9992 + w_sys_tmp9990);
	assign w_sys_tmp9992 = (r_run_copy6_j_277 * w_sys_tmp9969);
	assign w_sys_tmp9996 = (w_sys_tmp9997 + w_sys_tmp9999);
	assign w_sys_tmp9997 = (r_run_copy5_j_276 * w_sys_tmp9969);
	assign w_sys_tmp9999 = 32'sh00000040;
	assign w_sys_tmp10001 = (w_sys_tmp10002 + w_sys_tmp9999);
	assign w_sys_tmp10002 = (r_run_copy4_j_275 * w_sys_tmp9969);
	assign w_sys_tmp10006 = (w_sys_tmp10007 + w_sys_tmp10009);
	assign w_sys_tmp10007 = (r_run_copy3_j_274 * w_sys_tmp9969);
	assign w_sys_tmp10009 = 32'sh00000061;
	assign w_sys_tmp10010 = (w_sys_tmp10011 + w_sys_tmp10009);
	assign w_sys_tmp10011 = (r_run_copy2_j_273 * w_sys_tmp9969);
	assign w_sys_tmp10015 = (w_sys_tmp10016 + w_sys_tmp10018);
	assign w_sys_tmp10016 = (r_run_copy1_j_272 * w_sys_tmp9969);
	assign w_sys_tmp10018 = 32'sh00000060;
	assign w_sys_tmp10019 = w_sub21_result_dataout;
	assign w_sys_tmp10020 = (w_sys_tmp10021 + w_sys_tmp10018);
	assign w_sys_tmp10021 = (r_run_copy0_j_271 * w_sys_tmp9969);
	assign w_sys_tmp10024 = (r_run_copy0_j_271 + w_sys_intOne);
	assign w_sys_tmp10025 = (r_run_copy1_j_272 + w_sys_intOne);
	assign w_sys_tmp10026 = (r_run_copy2_j_273 + w_sys_intOne);
	assign w_sys_tmp10027 = (r_run_copy3_j_274 + w_sys_intOne);
	assign w_sys_tmp10028 = (r_run_copy4_j_275 + w_sys_intOne);
	assign w_sys_tmp10029 = (r_run_copy5_j_276 + w_sys_intOne);
	assign w_sys_tmp10030 = (r_run_copy6_j_277 + w_sys_intOne);
	assign w_sys_tmp10031 = (r_run_copy7_j_278 + w_sys_intOne);
	assign w_sys_tmp10032 = (r_run_copy8_j_279 + w_sys_intOne);
	assign w_sys_tmp10033 = (r_run_copy9_j_280 + w_sys_intOne);
	assign w_sys_tmp10034 = (r_run_copy10_j_281 + w_sys_intOne);
	assign w_sys_tmp10035 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp10462 = 32'sh00000060;
	assign w_sys_tmp10463 = ( !w_sys_tmp10464 );
	assign w_sys_tmp10464 = (w_sys_tmp10465 < r_run_j_37);
	assign w_sys_tmp10465 = 32'sh00000071;
	assign w_sys_tmp10468 = (w_sys_tmp10469 + w_sys_tmp10471);
	assign w_sys_tmp10469 = (r_run_j_37 * w_sys_tmp10470);
	assign w_sys_tmp10470 = 32'sh00000081;
	assign w_sys_tmp10471 = 32'sh00000021;
	assign w_sys_tmp10472 = w_sub14_result_dataout;
	assign w_sys_tmp10473 = (w_sys_tmp10474 + w_sys_tmp10471);
	assign w_sys_tmp10474 = (r_run_copy10_j_292 * w_sys_tmp10470);
	assign w_sys_tmp10478 = (w_sys_tmp10479 + w_sys_tmp10481);
	assign w_sys_tmp10479 = (r_run_copy9_j_291 * w_sys_tmp10470);
	assign w_sys_tmp10481 = 32'sh00000020;
	assign w_sys_tmp10482 = w_sub06_result_dataout;
	assign w_sys_tmp10483 = (w_sys_tmp10484 + w_sys_tmp10481);
	assign w_sys_tmp10484 = (r_run_copy8_j_290 * w_sys_tmp10470);
	assign w_sys_tmp10488 = (w_sys_tmp10489 + w_sys_tmp10491);
	assign w_sys_tmp10489 = (r_run_copy7_j_289 * w_sys_tmp10470);
	assign w_sys_tmp10491 = 32'sh00000041;
	assign w_sys_tmp10492 = (w_sys_tmp10493 + w_sys_tmp10491);
	assign w_sys_tmp10493 = (r_run_copy6_j_288 * w_sys_tmp10470);
	assign w_sys_tmp10497 = (w_sys_tmp10498 + w_sys_tmp10500);
	assign w_sys_tmp10498 = (r_run_copy5_j_287 * w_sys_tmp10470);
	assign w_sys_tmp10500 = 32'sh00000040;
	assign w_sys_tmp10502 = (w_sys_tmp10503 + w_sys_tmp10500);
	assign w_sys_tmp10503 = (r_run_copy4_j_286 * w_sys_tmp10470);
	assign w_sys_tmp10507 = (w_sys_tmp10508 + w_sys_tmp10510);
	assign w_sys_tmp10508 = (r_run_copy3_j_285 * w_sys_tmp10470);
	assign w_sys_tmp10510 = 32'sh00000061;
	assign w_sys_tmp10511 = (w_sys_tmp10512 + w_sys_tmp10510);
	assign w_sys_tmp10512 = (r_run_copy2_j_284 * w_sys_tmp10470);
	assign w_sys_tmp10516 = (w_sys_tmp10517 + w_sys_tmp10519);
	assign w_sys_tmp10517 = (r_run_copy1_j_283 * w_sys_tmp10470);
	assign w_sys_tmp10519 = 32'sh00000060;
	assign w_sys_tmp10520 = w_sub22_result_dataout;
	assign w_sys_tmp10521 = (w_sys_tmp10522 + w_sys_tmp10519);
	assign w_sys_tmp10522 = (r_run_copy0_j_282 * w_sys_tmp10470);
	assign w_sys_tmp10525 = (r_run_copy0_j_282 + w_sys_intOne);
	assign w_sys_tmp10526 = (r_run_copy1_j_283 + w_sys_intOne);
	assign w_sys_tmp10527 = (r_run_copy2_j_284 + w_sys_intOne);
	assign w_sys_tmp10528 = (r_run_copy3_j_285 + w_sys_intOne);
	assign w_sys_tmp10529 = (r_run_copy4_j_286 + w_sys_intOne);
	assign w_sys_tmp10530 = (r_run_copy5_j_287 + w_sys_intOne);
	assign w_sys_tmp10531 = (r_run_copy6_j_288 + w_sys_intOne);
	assign w_sys_tmp10532 = (r_run_copy7_j_289 + w_sys_intOne);
	assign w_sys_tmp10533 = (r_run_copy8_j_290 + w_sys_intOne);
	assign w_sys_tmp10534 = (r_run_copy9_j_291 + w_sys_intOne);
	assign w_sys_tmp10535 = (r_run_copy10_j_292 + w_sys_intOne);
	assign w_sys_tmp10536 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp10963 = 32'sh00000070;
	assign w_sys_tmp10964 = ( !w_sys_tmp10965 );
	assign w_sys_tmp10965 = (w_sys_tmp10966 < r_run_j_37);
	assign w_sys_tmp10966 = 32'sh00000081;
	assign w_sys_tmp10969 = (w_sys_tmp10970 + w_sys_tmp10972);
	assign w_sys_tmp10970 = (r_run_j_37 * w_sys_tmp10971);
	assign w_sys_tmp10971 = 32'sh00000081;
	assign w_sys_tmp10972 = 32'sh00000021;
	assign w_sys_tmp10973 = w_sub15_result_dataout;
	assign w_sys_tmp10974 = (w_sys_tmp10975 + w_sys_tmp10972);
	assign w_sys_tmp10975 = (r_run_copy10_j_303 * w_sys_tmp10971);
	assign w_sys_tmp10979 = (w_sys_tmp10980 + w_sys_tmp10982);
	assign w_sys_tmp10980 = (r_run_copy9_j_302 * w_sys_tmp10971);
	assign w_sys_tmp10982 = 32'sh00000020;
	assign w_sys_tmp10983 = w_sub07_result_dataout;
	assign w_sys_tmp10984 = (w_sys_tmp10985 + w_sys_tmp10982);
	assign w_sys_tmp10985 = (r_run_copy8_j_301 * w_sys_tmp10971);
	assign w_sys_tmp10989 = (w_sys_tmp10990 + w_sys_tmp10992);
	assign w_sys_tmp10990 = (r_run_copy7_j_300 * w_sys_tmp10971);
	assign w_sys_tmp10992 = 32'sh00000041;
	assign w_sys_tmp10993 = (w_sys_tmp10994 + w_sys_tmp10992);
	assign w_sys_tmp10994 = (r_run_copy6_j_299 * w_sys_tmp10971);
	assign w_sys_tmp10998 = (w_sys_tmp10999 + w_sys_tmp11001);
	assign w_sys_tmp10999 = (r_run_copy5_j_298 * w_sys_tmp10971);
	assign w_sys_tmp11001 = 32'sh00000040;
	assign w_sys_tmp11003 = (w_sys_tmp11004 + w_sys_tmp11001);
	assign w_sys_tmp11004 = (r_run_copy4_j_297 * w_sys_tmp10971);
	assign w_sys_tmp11008 = (w_sys_tmp11009 + w_sys_tmp11011);
	assign w_sys_tmp11009 = (r_run_copy3_j_296 * w_sys_tmp10971);
	assign w_sys_tmp11011 = 32'sh00000061;
	assign w_sys_tmp11012 = (w_sys_tmp11013 + w_sys_tmp11011);
	assign w_sys_tmp11013 = (r_run_copy2_j_295 * w_sys_tmp10971);
	assign w_sys_tmp11017 = (w_sys_tmp11018 + w_sys_tmp11020);
	assign w_sys_tmp11018 = (r_run_copy1_j_294 * w_sys_tmp10971);
	assign w_sys_tmp11020 = 32'sh00000060;
	assign w_sys_tmp11021 = w_sub16_result_dataout;
	assign w_sys_tmp11022 = (w_sys_tmp11023 + w_sys_tmp11020);
	assign w_sys_tmp11023 = (r_run_copy0_j_293 * w_sys_tmp10971);
	assign w_sys_tmp11026 = (r_run_copy0_j_293 + w_sys_intOne);
	assign w_sys_tmp11027 = (r_run_copy1_j_294 + w_sys_intOne);
	assign w_sys_tmp11028 = (r_run_copy2_j_295 + w_sys_intOne);
	assign w_sys_tmp11029 = (r_run_copy3_j_296 + w_sys_intOne);
	assign w_sys_tmp11030 = (r_run_copy4_j_297 + w_sys_intOne);
	assign w_sys_tmp11031 = (r_run_copy5_j_298 + w_sys_intOne);
	assign w_sys_tmp11032 = (r_run_copy6_j_299 + w_sys_intOne);
	assign w_sys_tmp11033 = (r_run_copy7_j_300 + w_sys_intOne);
	assign w_sys_tmp11034 = (r_run_copy8_j_301 + w_sys_intOne);
	assign w_sys_tmp11035 = (r_run_copy9_j_302 + w_sys_intOne);
	assign w_sys_tmp11036 = (r_run_copy10_j_303 + w_sys_intOne);
	assign w_sys_tmp11037 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp11452 = 32'sh00000002;
	assign w_sys_tmp11453 = ( !w_sys_tmp11454 );
	assign w_sys_tmp11454 = (w_sys_tmp11455 < r_run_k_36);
	assign w_sys_tmp11455 = 32'sh00000020;
	assign w_sys_tmp11456 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp11457 = 32'sh00000002;
	assign w_sys_tmp11458 = ( !w_sys_tmp11459 );
	assign w_sys_tmp11459 = (w_sys_tmp11460 < r_run_j_37);
	assign w_sys_tmp11460 = 32'sh00000010;
	assign w_sys_tmp11463 = (w_sys_tmp11464 + r_run_k_36);
	assign w_sys_tmp11464 = (r_run_j_37 * w_sys_tmp11465);
	assign w_sys_tmp11465 = 32'sh00000081;
	assign w_sys_tmp11466 = w_sub00_result_dataout;
	assign w_sys_tmp11467 = (w_sys_tmp11468 + r_run_k_36);
	assign w_sys_tmp11468 = (r_run_copy0_j_304 * w_sys_tmp11465);
	assign w_sys_tmp11470 = (r_run_copy0_j_304 + w_sys_intOne);
	assign w_sys_tmp11471 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp11532 = 32'sh00000011;
	assign w_sys_tmp11533 = ( !w_sys_tmp11534 );
	assign w_sys_tmp11534 = (w_sys_tmp11535 < r_run_j_37);
	assign w_sys_tmp11535 = 32'sh00000020;
	assign w_sys_tmp11537 = (r_run_j_37 - w_sys_tmp11538);
	assign w_sys_tmp11538 = 32'sh0000000f;
	assign w_sys_tmp11540 = (w_sys_tmp11541 + r_run_k_36);
	assign w_sys_tmp11541 = (r_run_copy1_j_306 * w_sys_tmp11542);
	assign w_sys_tmp11542 = 32'sh00000081;
	assign w_sys_tmp11543 = w_sub01_result_dataout;
	assign w_sys_tmp11544 = (w_sys_tmp11545 + r_run_k_36);
	assign w_sys_tmp11545 = (r_run_copy0_j_305 * w_sys_tmp11542);
	assign w_sys_tmp11547 = (r_run_copy0_j_305 + w_sys_intOne);
	assign w_sys_tmp11548 = (r_run_copy1_j_306 + w_sys_intOne);
	assign w_sys_tmp11549 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp11628 = 32'sh00000021;
	assign w_sys_tmp11629 = ( !w_sys_tmp11630 );
	assign w_sys_tmp11630 = (w_sys_tmp11631 < r_run_j_37);
	assign w_sys_tmp11631 = 32'sh00000030;
	assign w_sys_tmp11633 = (r_run_j_37 - w_sys_tmp11634);
	assign w_sys_tmp11634 = 32'sh0000001f;
	assign w_sys_tmp11636 = (w_sys_tmp11637 + r_run_k_36);
	assign w_sys_tmp11637 = (r_run_copy1_j_308 * w_sys_tmp11638);
	assign w_sys_tmp11638 = 32'sh00000081;
	assign w_sys_tmp11639 = w_sub02_result_dataout;
	assign w_sys_tmp11640 = (w_sys_tmp11641 + r_run_k_36);
	assign w_sys_tmp11641 = (r_run_copy0_j_307 * w_sys_tmp11638);
	assign w_sys_tmp11643 = (r_run_copy0_j_307 + w_sys_intOne);
	assign w_sys_tmp11644 = (r_run_copy1_j_308 + w_sys_intOne);
	assign w_sys_tmp11645 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp11724 = 32'sh00000031;
	assign w_sys_tmp11725 = ( !w_sys_tmp11726 );
	assign w_sys_tmp11726 = (w_sys_tmp11727 < r_run_j_37);
	assign w_sys_tmp11727 = 32'sh00000040;
	assign w_sys_tmp11729 = (r_run_j_37 - w_sys_tmp11730);
	assign w_sys_tmp11730 = 32'sh0000002f;
	assign w_sys_tmp11732 = (w_sys_tmp11733 + r_run_k_36);
	assign w_sys_tmp11733 = (r_run_copy1_j_310 * w_sys_tmp11734);
	assign w_sys_tmp11734 = 32'sh00000081;
	assign w_sys_tmp11735 = w_sub03_result_dataout;
	assign w_sys_tmp11736 = (w_sys_tmp11737 + r_run_k_36);
	assign w_sys_tmp11737 = (r_run_copy0_j_309 * w_sys_tmp11734);
	assign w_sys_tmp11739 = (r_run_copy0_j_309 + w_sys_intOne);
	assign w_sys_tmp11740 = (r_run_copy1_j_310 + w_sys_intOne);
	assign w_sys_tmp11741 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp11820 = 32'sh00000041;
	assign w_sys_tmp11821 = ( !w_sys_tmp11822 );
	assign w_sys_tmp11822 = (w_sys_tmp11823 < r_run_j_37);
	assign w_sys_tmp11823 = 32'sh00000050;
	assign w_sys_tmp11825 = (r_run_j_37 - w_sys_tmp11826);
	assign w_sys_tmp11826 = 32'sh0000003f;
	assign w_sys_tmp11828 = (w_sys_tmp11829 + r_run_k_36);
	assign w_sys_tmp11829 = (r_run_copy1_j_312 * w_sys_tmp11830);
	assign w_sys_tmp11830 = 32'sh00000081;
	assign w_sys_tmp11831 = w_sub04_result_dataout;
	assign w_sys_tmp11832 = (w_sys_tmp11833 + r_run_k_36);
	assign w_sys_tmp11833 = (r_run_copy0_j_311 * w_sys_tmp11830);
	assign w_sys_tmp11835 = (r_run_copy0_j_311 + w_sys_intOne);
	assign w_sys_tmp11836 = (r_run_copy1_j_312 + w_sys_intOne);
	assign w_sys_tmp11837 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp11916 = 32'sh00000051;
	assign w_sys_tmp11917 = ( !w_sys_tmp11918 );
	assign w_sys_tmp11918 = (w_sys_tmp11919 < r_run_j_37);
	assign w_sys_tmp11919 = 32'sh00000060;
	assign w_sys_tmp11921 = (r_run_j_37 - w_sys_tmp11922);
	assign w_sys_tmp11922 = 32'sh0000004f;
	assign w_sys_tmp11924 = (w_sys_tmp11925 + r_run_k_36);
	assign w_sys_tmp11925 = (r_run_copy1_j_314 * w_sys_tmp11926);
	assign w_sys_tmp11926 = 32'sh00000081;
	assign w_sys_tmp11927 = w_sub05_result_dataout;
	assign w_sys_tmp11928 = (w_sys_tmp11929 + r_run_k_36);
	assign w_sys_tmp11929 = (r_run_copy0_j_313 * w_sys_tmp11926);
	assign w_sys_tmp11931 = (r_run_copy0_j_313 + w_sys_intOne);
	assign w_sys_tmp11932 = (r_run_copy1_j_314 + w_sys_intOne);
	assign w_sys_tmp11933 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12012 = 32'sh00000061;
	assign w_sys_tmp12013 = ( !w_sys_tmp12014 );
	assign w_sys_tmp12014 = (w_sys_tmp12015 < r_run_j_37);
	assign w_sys_tmp12015 = 32'sh00000070;
	assign w_sys_tmp12017 = (r_run_j_37 - w_sys_tmp12018);
	assign w_sys_tmp12018 = 32'sh0000005f;
	assign w_sys_tmp12020 = (w_sys_tmp12021 + r_run_k_36);
	assign w_sys_tmp12021 = (r_run_copy1_j_316 * w_sys_tmp12022);
	assign w_sys_tmp12022 = 32'sh00000081;
	assign w_sys_tmp12023 = w_sub06_result_dataout;
	assign w_sys_tmp12024 = (w_sys_tmp12025 + r_run_k_36);
	assign w_sys_tmp12025 = (r_run_copy0_j_315 * w_sys_tmp12022);
	assign w_sys_tmp12027 = (r_run_copy0_j_315 + w_sys_intOne);
	assign w_sys_tmp12028 = (r_run_copy1_j_316 + w_sys_intOne);
	assign w_sys_tmp12029 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12108 = 32'sh00000071;
	assign w_sys_tmp12109 = ( !w_sys_tmp12110 );
	assign w_sys_tmp12110 = (w_sys_tmp12111 < r_run_j_37);
	assign w_sys_tmp12111 = 32'sh00000080;
	assign w_sys_tmp12113 = (r_run_j_37 - w_sys_tmp12114);
	assign w_sys_tmp12114 = 32'sh0000006f;
	assign w_sys_tmp12116 = (w_sys_tmp12117 + r_run_k_36);
	assign w_sys_tmp12117 = (r_run_copy1_j_318 * w_sys_tmp12118);
	assign w_sys_tmp12118 = 32'sh00000081;
	assign w_sys_tmp12119 = w_sub07_result_dataout;
	assign w_sys_tmp12120 = (w_sys_tmp12121 + r_run_k_36);
	assign w_sys_tmp12121 = (r_run_copy0_j_317 * w_sys_tmp12118);
	assign w_sys_tmp12123 = (r_run_copy0_j_317 + w_sys_intOne);
	assign w_sys_tmp12124 = (r_run_copy1_j_318 + w_sys_intOne);
	assign w_sys_tmp12125 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12204 = 32'sh00000021;
	assign w_sys_tmp12205 = ( !w_sys_tmp12206 );
	assign w_sys_tmp12206 = (w_sys_tmp12207 < r_run_k_36);
	assign w_sys_tmp12207 = 32'sh00000040;
	assign w_sys_tmp12208 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp12209 = 32'sh00000002;
	assign w_sys_tmp12210 = ( !w_sys_tmp12211 );
	assign w_sys_tmp12211 = (w_sys_tmp12212 < r_run_j_37);
	assign w_sys_tmp12212 = 32'sh00000010;
	assign w_sys_tmp12215 = (w_sys_tmp12216 + r_run_k_36);
	assign w_sys_tmp12216 = (r_run_j_37 * w_sys_tmp12217);
	assign w_sys_tmp12217 = 32'sh00000081;
	assign w_sys_tmp12218 = w_sub08_result_dataout;
	assign w_sys_tmp12219 = (w_sys_tmp12220 + r_run_k_36);
	assign w_sys_tmp12220 = (r_run_copy0_j_319 * w_sys_tmp12217);
	assign w_sys_tmp12222 = (r_run_copy0_j_319 + w_sys_intOne);
	assign w_sys_tmp12223 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12284 = 32'sh00000011;
	assign w_sys_tmp12285 = ( !w_sys_tmp12286 );
	assign w_sys_tmp12286 = (w_sys_tmp12287 < r_run_j_37);
	assign w_sys_tmp12287 = 32'sh00000020;
	assign w_sys_tmp12289 = (r_run_j_37 - w_sys_tmp12290);
	assign w_sys_tmp12290 = 32'sh0000000f;
	assign w_sys_tmp12292 = (w_sys_tmp12293 + r_run_k_36);
	assign w_sys_tmp12293 = (r_run_copy1_j_321 * w_sys_tmp12294);
	assign w_sys_tmp12294 = 32'sh00000081;
	assign w_sys_tmp12295 = w_sub09_result_dataout;
	assign w_sys_tmp12296 = (w_sys_tmp12297 + r_run_k_36);
	assign w_sys_tmp12297 = (r_run_copy0_j_320 * w_sys_tmp12294);
	assign w_sys_tmp12299 = (r_run_copy0_j_320 + w_sys_intOne);
	assign w_sys_tmp12300 = (r_run_copy1_j_321 + w_sys_intOne);
	assign w_sys_tmp12301 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12380 = 32'sh00000021;
	assign w_sys_tmp12381 = ( !w_sys_tmp12382 );
	assign w_sys_tmp12382 = (w_sys_tmp12383 < r_run_j_37);
	assign w_sys_tmp12383 = 32'sh00000030;
	assign w_sys_tmp12385 = (r_run_j_37 - w_sys_tmp12386);
	assign w_sys_tmp12386 = 32'sh0000001f;
	assign w_sys_tmp12388 = (w_sys_tmp12389 + r_run_k_36);
	assign w_sys_tmp12389 = (r_run_copy1_j_323 * w_sys_tmp12390);
	assign w_sys_tmp12390 = 32'sh00000081;
	assign w_sys_tmp12391 = w_sub10_result_dataout;
	assign w_sys_tmp12392 = (w_sys_tmp12393 + r_run_k_36);
	assign w_sys_tmp12393 = (r_run_copy0_j_322 * w_sys_tmp12390);
	assign w_sys_tmp12395 = (r_run_copy0_j_322 + w_sys_intOne);
	assign w_sys_tmp12396 = (r_run_copy1_j_323 + w_sys_intOne);
	assign w_sys_tmp12397 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12476 = 32'sh00000031;
	assign w_sys_tmp12477 = ( !w_sys_tmp12478 );
	assign w_sys_tmp12478 = (w_sys_tmp12479 < r_run_j_37);
	assign w_sys_tmp12479 = 32'sh00000040;
	assign w_sys_tmp12481 = (r_run_j_37 - w_sys_tmp12482);
	assign w_sys_tmp12482 = 32'sh0000002f;
	assign w_sys_tmp12484 = (w_sys_tmp12485 + r_run_k_36);
	assign w_sys_tmp12485 = (r_run_copy1_j_325 * w_sys_tmp12486);
	assign w_sys_tmp12486 = 32'sh00000081;
	assign w_sys_tmp12487 = w_sub11_result_dataout;
	assign w_sys_tmp12488 = (w_sys_tmp12489 + r_run_k_36);
	assign w_sys_tmp12489 = (r_run_copy0_j_324 * w_sys_tmp12486);
	assign w_sys_tmp12491 = (r_run_copy0_j_324 + w_sys_intOne);
	assign w_sys_tmp12492 = (r_run_copy1_j_325 + w_sys_intOne);
	assign w_sys_tmp12493 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12572 = 32'sh00000041;
	assign w_sys_tmp12573 = ( !w_sys_tmp12574 );
	assign w_sys_tmp12574 = (w_sys_tmp12575 < r_run_j_37);
	assign w_sys_tmp12575 = 32'sh00000050;
	assign w_sys_tmp12577 = (r_run_j_37 - w_sys_tmp12578);
	assign w_sys_tmp12578 = 32'sh0000003f;
	assign w_sys_tmp12580 = (w_sys_tmp12581 + r_run_k_36);
	assign w_sys_tmp12581 = (r_run_copy1_j_327 * w_sys_tmp12582);
	assign w_sys_tmp12582 = 32'sh00000081;
	assign w_sys_tmp12583 = w_sub12_result_dataout;
	assign w_sys_tmp12584 = (w_sys_tmp12585 + r_run_k_36);
	assign w_sys_tmp12585 = (r_run_copy0_j_326 * w_sys_tmp12582);
	assign w_sys_tmp12587 = (r_run_copy0_j_326 + w_sys_intOne);
	assign w_sys_tmp12588 = (r_run_copy1_j_327 + w_sys_intOne);
	assign w_sys_tmp12589 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12668 = 32'sh00000051;
	assign w_sys_tmp12669 = ( !w_sys_tmp12670 );
	assign w_sys_tmp12670 = (w_sys_tmp12671 < r_run_j_37);
	assign w_sys_tmp12671 = 32'sh00000060;
	assign w_sys_tmp12673 = (r_run_j_37 - w_sys_tmp12674);
	assign w_sys_tmp12674 = 32'sh0000004f;
	assign w_sys_tmp12676 = (w_sys_tmp12677 + r_run_k_36);
	assign w_sys_tmp12677 = (r_run_copy1_j_329 * w_sys_tmp12678);
	assign w_sys_tmp12678 = 32'sh00000081;
	assign w_sys_tmp12679 = w_sub13_result_dataout;
	assign w_sys_tmp12680 = (w_sys_tmp12681 + r_run_k_36);
	assign w_sys_tmp12681 = (r_run_copy0_j_328 * w_sys_tmp12678);
	assign w_sys_tmp12683 = (r_run_copy0_j_328 + w_sys_intOne);
	assign w_sys_tmp12684 = (r_run_copy1_j_329 + w_sys_intOne);
	assign w_sys_tmp12685 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12764 = 32'sh00000061;
	assign w_sys_tmp12765 = ( !w_sys_tmp12766 );
	assign w_sys_tmp12766 = (w_sys_tmp12767 < r_run_j_37);
	assign w_sys_tmp12767 = 32'sh00000070;
	assign w_sys_tmp12769 = (r_run_j_37 - w_sys_tmp12770);
	assign w_sys_tmp12770 = 32'sh0000005f;
	assign w_sys_tmp12772 = (w_sys_tmp12773 + r_run_k_36);
	assign w_sys_tmp12773 = (r_run_copy1_j_331 * w_sys_tmp12774);
	assign w_sys_tmp12774 = 32'sh00000081;
	assign w_sys_tmp12775 = w_sub14_result_dataout;
	assign w_sys_tmp12776 = (w_sys_tmp12777 + r_run_k_36);
	assign w_sys_tmp12777 = (r_run_copy0_j_330 * w_sys_tmp12774);
	assign w_sys_tmp12779 = (r_run_copy0_j_330 + w_sys_intOne);
	assign w_sys_tmp12780 = (r_run_copy1_j_331 + w_sys_intOne);
	assign w_sys_tmp12781 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12860 = 32'sh00000071;
	assign w_sys_tmp12861 = ( !w_sys_tmp12862 );
	assign w_sys_tmp12862 = (w_sys_tmp12863 < r_run_j_37);
	assign w_sys_tmp12863 = 32'sh00000080;
	assign w_sys_tmp12865 = (r_run_j_37 - w_sys_tmp12866);
	assign w_sys_tmp12866 = 32'sh0000006f;
	assign w_sys_tmp12868 = (w_sys_tmp12869 + r_run_k_36);
	assign w_sys_tmp12869 = (r_run_copy1_j_333 * w_sys_tmp12870);
	assign w_sys_tmp12870 = 32'sh00000081;
	assign w_sys_tmp12871 = w_sub15_result_dataout;
	assign w_sys_tmp12872 = (w_sys_tmp12873 + r_run_k_36);
	assign w_sys_tmp12873 = (r_run_copy0_j_332 * w_sys_tmp12870);
	assign w_sys_tmp12875 = (r_run_copy0_j_332 + w_sys_intOne);
	assign w_sys_tmp12876 = (r_run_copy1_j_333 + w_sys_intOne);
	assign w_sys_tmp12877 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp12956 = 32'sh00000041;
	assign w_sys_tmp12957 = ( !w_sys_tmp12958 );
	assign w_sys_tmp12958 = (w_sys_tmp12959 < r_run_k_36);
	assign w_sys_tmp12959 = 32'sh00000060;
	assign w_sys_tmp12960 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp12961 = 32'sh00000002;
	assign w_sys_tmp12962 = ( !w_sys_tmp12963 );
	assign w_sys_tmp12963 = (w_sys_tmp12964 < r_run_j_37);
	assign w_sys_tmp12964 = 32'sh00000010;
	assign w_sys_tmp12967 = (w_sys_tmp12968 + r_run_k_36);
	assign w_sys_tmp12968 = (r_run_j_37 * w_sys_tmp12969);
	assign w_sys_tmp12969 = 32'sh00000081;
	assign w_sys_tmp12970 = w_sub16_result_dataout;
	assign w_sys_tmp12971 = (w_sys_tmp12972 + r_run_k_36);
	assign w_sys_tmp12972 = (r_run_copy0_j_334 * w_sys_tmp12969);
	assign w_sys_tmp12974 = (r_run_copy0_j_334 + w_sys_intOne);
	assign w_sys_tmp12975 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13036 = 32'sh00000011;
	assign w_sys_tmp13037 = ( !w_sys_tmp13038 );
	assign w_sys_tmp13038 = (w_sys_tmp13039 < r_run_j_37);
	assign w_sys_tmp13039 = 32'sh00000020;
	assign w_sys_tmp13041 = (r_run_j_37 - w_sys_tmp13042);
	assign w_sys_tmp13042 = 32'sh0000000f;
	assign w_sys_tmp13044 = (w_sys_tmp13045 + r_run_k_36);
	assign w_sys_tmp13045 = (r_run_copy1_j_336 * w_sys_tmp13046);
	assign w_sys_tmp13046 = 32'sh00000081;
	assign w_sys_tmp13047 = w_sub17_result_dataout;
	assign w_sys_tmp13048 = (w_sys_tmp13049 + r_run_k_36);
	assign w_sys_tmp13049 = (r_run_copy0_j_335 * w_sys_tmp13046);
	assign w_sys_tmp13051 = (r_run_copy0_j_335 + w_sys_intOne);
	assign w_sys_tmp13052 = (r_run_copy1_j_336 + w_sys_intOne);
	assign w_sys_tmp13053 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13132 = 32'sh00000021;
	assign w_sys_tmp13133 = ( !w_sys_tmp13134 );
	assign w_sys_tmp13134 = (w_sys_tmp13135 < r_run_j_37);
	assign w_sys_tmp13135 = 32'sh00000030;
	assign w_sys_tmp13137 = (r_run_j_37 - w_sys_tmp13138);
	assign w_sys_tmp13138 = 32'sh0000001f;
	assign w_sys_tmp13140 = (w_sys_tmp13141 + r_run_k_36);
	assign w_sys_tmp13141 = (r_run_copy1_j_338 * w_sys_tmp13142);
	assign w_sys_tmp13142 = 32'sh00000081;
	assign w_sys_tmp13143 = w_sub18_result_dataout;
	assign w_sys_tmp13144 = (w_sys_tmp13145 + r_run_k_36);
	assign w_sys_tmp13145 = (r_run_copy0_j_337 * w_sys_tmp13142);
	assign w_sys_tmp13147 = (r_run_copy0_j_337 + w_sys_intOne);
	assign w_sys_tmp13148 = (r_run_copy1_j_338 + w_sys_intOne);
	assign w_sys_tmp13149 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13228 = 32'sh00000031;
	assign w_sys_tmp13229 = ( !w_sys_tmp13230 );
	assign w_sys_tmp13230 = (w_sys_tmp13231 < r_run_j_37);
	assign w_sys_tmp13231 = 32'sh00000040;
	assign w_sys_tmp13233 = (r_run_j_37 - w_sys_tmp13234);
	assign w_sys_tmp13234 = 32'sh0000002f;
	assign w_sys_tmp13236 = (w_sys_tmp13237 + r_run_k_36);
	assign w_sys_tmp13237 = (r_run_copy1_j_340 * w_sys_tmp13238);
	assign w_sys_tmp13238 = 32'sh00000081;
	assign w_sys_tmp13239 = w_sub19_result_dataout;
	assign w_sys_tmp13240 = (w_sys_tmp13241 + r_run_k_36);
	assign w_sys_tmp13241 = (r_run_copy0_j_339 * w_sys_tmp13238);
	assign w_sys_tmp13243 = (r_run_copy0_j_339 + w_sys_intOne);
	assign w_sys_tmp13244 = (r_run_copy1_j_340 + w_sys_intOne);
	assign w_sys_tmp13245 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13324 = 32'sh00000041;
	assign w_sys_tmp13325 = ( !w_sys_tmp13326 );
	assign w_sys_tmp13326 = (w_sys_tmp13327 < r_run_j_37);
	assign w_sys_tmp13327 = 32'sh00000050;
	assign w_sys_tmp13329 = (r_run_j_37 - w_sys_tmp13330);
	assign w_sys_tmp13330 = 32'sh0000003f;
	assign w_sys_tmp13332 = (w_sys_tmp13333 + r_run_k_36);
	assign w_sys_tmp13333 = (r_run_copy1_j_342 * w_sys_tmp13334);
	assign w_sys_tmp13334 = 32'sh00000081;
	assign w_sys_tmp13335 = w_sub20_result_dataout;
	assign w_sys_tmp13336 = (w_sys_tmp13337 + r_run_k_36);
	assign w_sys_tmp13337 = (r_run_copy0_j_341 * w_sys_tmp13334);
	assign w_sys_tmp13339 = (r_run_copy0_j_341 + w_sys_intOne);
	assign w_sys_tmp13340 = (r_run_copy1_j_342 + w_sys_intOne);
	assign w_sys_tmp13341 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13420 = 32'sh00000051;
	assign w_sys_tmp13421 = ( !w_sys_tmp13422 );
	assign w_sys_tmp13422 = (w_sys_tmp13423 < r_run_j_37);
	assign w_sys_tmp13423 = 32'sh00000060;
	assign w_sys_tmp13425 = (r_run_j_37 - w_sys_tmp13426);
	assign w_sys_tmp13426 = 32'sh0000004f;
	assign w_sys_tmp13428 = (w_sys_tmp13429 + r_run_k_36);
	assign w_sys_tmp13429 = (r_run_copy1_j_344 * w_sys_tmp13430);
	assign w_sys_tmp13430 = 32'sh00000081;
	assign w_sys_tmp13431 = w_sub21_result_dataout;
	assign w_sys_tmp13432 = (w_sys_tmp13433 + r_run_k_36);
	assign w_sys_tmp13433 = (r_run_copy0_j_343 * w_sys_tmp13430);
	assign w_sys_tmp13435 = (r_run_copy0_j_343 + w_sys_intOne);
	assign w_sys_tmp13436 = (r_run_copy1_j_344 + w_sys_intOne);
	assign w_sys_tmp13437 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13516 = 32'sh00000061;
	assign w_sys_tmp13517 = ( !w_sys_tmp13518 );
	assign w_sys_tmp13518 = (w_sys_tmp13519 < r_run_j_37);
	assign w_sys_tmp13519 = 32'sh00000070;
	assign w_sys_tmp13521 = (r_run_j_37 - w_sys_tmp13522);
	assign w_sys_tmp13522 = 32'sh0000005f;
	assign w_sys_tmp13524 = (w_sys_tmp13525 + r_run_k_36);
	assign w_sys_tmp13525 = (r_run_copy1_j_346 * w_sys_tmp13526);
	assign w_sys_tmp13526 = 32'sh00000081;
	assign w_sys_tmp13527 = w_sub22_result_dataout;
	assign w_sys_tmp13528 = (w_sys_tmp13529 + r_run_k_36);
	assign w_sys_tmp13529 = (r_run_copy0_j_345 * w_sys_tmp13526);
	assign w_sys_tmp13531 = (r_run_copy0_j_345 + w_sys_intOne);
	assign w_sys_tmp13532 = (r_run_copy1_j_346 + w_sys_intOne);
	assign w_sys_tmp13533 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13612 = 32'sh00000071;
	assign w_sys_tmp13613 = ( !w_sys_tmp13614 );
	assign w_sys_tmp13614 = (w_sys_tmp13615 < r_run_j_37);
	assign w_sys_tmp13615 = 32'sh00000080;
	assign w_sys_tmp13617 = (r_run_j_37 - w_sys_tmp13618);
	assign w_sys_tmp13618 = 32'sh0000006f;
	assign w_sys_tmp13620 = (w_sys_tmp13621 + r_run_k_36);
	assign w_sys_tmp13621 = (r_run_copy1_j_348 * w_sys_tmp13622);
	assign w_sys_tmp13622 = 32'sh00000081;
	assign w_sys_tmp13623 = w_sub23_result_dataout;
	assign w_sys_tmp13624 = (w_sys_tmp13625 + r_run_k_36);
	assign w_sys_tmp13625 = (r_run_copy0_j_347 * w_sys_tmp13622);
	assign w_sys_tmp13627 = (r_run_copy0_j_347 + w_sys_intOne);
	assign w_sys_tmp13628 = (r_run_copy1_j_348 + w_sys_intOne);
	assign w_sys_tmp13629 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13708 = 32'sh00000061;
	assign w_sys_tmp13709 = ( !w_sys_tmp13710 );
	assign w_sys_tmp13710 = (w_sys_tmp13711 < r_run_k_36);
	assign w_sys_tmp13711 = 32'sh00000080;
	assign w_sys_tmp13712 = (r_run_k_36 + w_sys_intOne);
	assign w_sys_tmp13713 = 32'sh00000002;
	assign w_sys_tmp13714 = ( !w_sys_tmp13715 );
	assign w_sys_tmp13715 = (w_sys_tmp13716 < r_run_j_37);
	assign w_sys_tmp13716 = 32'sh00000010;
	assign w_sys_tmp13719 = (w_sys_tmp13720 + r_run_k_36);
	assign w_sys_tmp13720 = (r_run_j_37 * w_sys_tmp13721);
	assign w_sys_tmp13721 = 32'sh00000081;
	assign w_sys_tmp13722 = w_sub24_result_dataout;
	assign w_sys_tmp13723 = (w_sys_tmp13724 + r_run_k_36);
	assign w_sys_tmp13724 = (r_run_copy0_j_349 * w_sys_tmp13721);
	assign w_sys_tmp13726 = (r_run_copy0_j_349 + w_sys_intOne);
	assign w_sys_tmp13727 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13788 = 32'sh00000011;
	assign w_sys_tmp13789 = ( !w_sys_tmp13790 );
	assign w_sys_tmp13790 = (w_sys_tmp13791 < r_run_j_37);
	assign w_sys_tmp13791 = 32'sh00000020;
	assign w_sys_tmp13793 = (r_run_j_37 - w_sys_tmp13794);
	assign w_sys_tmp13794 = 32'sh0000000f;
	assign w_sys_tmp13796 = (w_sys_tmp13797 + r_run_k_36);
	assign w_sys_tmp13797 = (r_run_copy1_j_351 * w_sys_tmp13798);
	assign w_sys_tmp13798 = 32'sh00000081;
	assign w_sys_tmp13799 = w_sub25_result_dataout;
	assign w_sys_tmp13800 = (w_sys_tmp13801 + r_run_k_36);
	assign w_sys_tmp13801 = (r_run_copy0_j_350 * w_sys_tmp13798);
	assign w_sys_tmp13803 = (r_run_copy0_j_350 + w_sys_intOne);
	assign w_sys_tmp13804 = (r_run_copy1_j_351 + w_sys_intOne);
	assign w_sys_tmp13805 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13884 = 32'sh00000021;
	assign w_sys_tmp13885 = ( !w_sys_tmp13886 );
	assign w_sys_tmp13886 = (w_sys_tmp13887 < r_run_j_37);
	assign w_sys_tmp13887 = 32'sh00000030;
	assign w_sys_tmp13889 = (r_run_j_37 - w_sys_tmp13890);
	assign w_sys_tmp13890 = 32'sh0000001f;
	assign w_sys_tmp13892 = (w_sys_tmp13893 + r_run_k_36);
	assign w_sys_tmp13893 = (r_run_copy1_j_353 * w_sys_tmp13894);
	assign w_sys_tmp13894 = 32'sh00000081;
	assign w_sys_tmp13895 = w_sub26_result_dataout;
	assign w_sys_tmp13896 = (w_sys_tmp13897 + r_run_k_36);
	assign w_sys_tmp13897 = (r_run_copy0_j_352 * w_sys_tmp13894);
	assign w_sys_tmp13899 = (r_run_copy0_j_352 + w_sys_intOne);
	assign w_sys_tmp13900 = (r_run_copy1_j_353 + w_sys_intOne);
	assign w_sys_tmp13901 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp13980 = 32'sh00000031;
	assign w_sys_tmp13981 = ( !w_sys_tmp13982 );
	assign w_sys_tmp13982 = (w_sys_tmp13983 < r_run_j_37);
	assign w_sys_tmp13983 = 32'sh00000040;
	assign w_sys_tmp13985 = (r_run_j_37 - w_sys_tmp13986);
	assign w_sys_tmp13986 = 32'sh0000002f;
	assign w_sys_tmp13988 = (w_sys_tmp13989 + r_run_k_36);
	assign w_sys_tmp13989 = (r_run_copy1_j_355 * w_sys_tmp13990);
	assign w_sys_tmp13990 = 32'sh00000081;
	assign w_sys_tmp13991 = w_sub27_result_dataout;
	assign w_sys_tmp13992 = (w_sys_tmp13993 + r_run_k_36);
	assign w_sys_tmp13993 = (r_run_copy0_j_354 * w_sys_tmp13990);
	assign w_sys_tmp13995 = (r_run_copy0_j_354 + w_sys_intOne);
	assign w_sys_tmp13996 = (r_run_copy1_j_355 + w_sys_intOne);
	assign w_sys_tmp13997 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp14076 = 32'sh00000041;
	assign w_sys_tmp14077 = ( !w_sys_tmp14078 );
	assign w_sys_tmp14078 = (w_sys_tmp14079 < r_run_j_37);
	assign w_sys_tmp14079 = 32'sh00000050;
	assign w_sys_tmp14081 = (r_run_j_37 - w_sys_tmp14082);
	assign w_sys_tmp14082 = 32'sh0000003f;
	assign w_sys_tmp14084 = (w_sys_tmp14085 + r_run_k_36);
	assign w_sys_tmp14085 = (r_run_copy1_j_357 * w_sys_tmp14086);
	assign w_sys_tmp14086 = 32'sh00000081;
	assign w_sys_tmp14087 = w_sub28_result_dataout;
	assign w_sys_tmp14088 = (w_sys_tmp14089 + r_run_k_36);
	assign w_sys_tmp14089 = (r_run_copy0_j_356 * w_sys_tmp14086);
	assign w_sys_tmp14091 = (r_run_copy0_j_356 + w_sys_intOne);
	assign w_sys_tmp14092 = (r_run_copy1_j_357 + w_sys_intOne);
	assign w_sys_tmp14093 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp14172 = 32'sh00000051;
	assign w_sys_tmp14173 = ( !w_sys_tmp14174 );
	assign w_sys_tmp14174 = (w_sys_tmp14175 < r_run_j_37);
	assign w_sys_tmp14175 = 32'sh00000060;
	assign w_sys_tmp14177 = (r_run_j_37 - w_sys_tmp14178);
	assign w_sys_tmp14178 = 32'sh0000004f;
	assign w_sys_tmp14180 = (w_sys_tmp14181 + r_run_k_36);
	assign w_sys_tmp14181 = (r_run_copy1_j_359 * w_sys_tmp14182);
	assign w_sys_tmp14182 = 32'sh00000081;
	assign w_sys_tmp14183 = w_sub29_result_dataout;
	assign w_sys_tmp14184 = (w_sys_tmp14185 + r_run_k_36);
	assign w_sys_tmp14185 = (r_run_copy0_j_358 * w_sys_tmp14182);
	assign w_sys_tmp14187 = (r_run_copy0_j_358 + w_sys_intOne);
	assign w_sys_tmp14188 = (r_run_copy1_j_359 + w_sys_intOne);
	assign w_sys_tmp14189 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp14268 = 32'sh00000061;
	assign w_sys_tmp14269 = ( !w_sys_tmp14270 );
	assign w_sys_tmp14270 = (w_sys_tmp14271 < r_run_j_37);
	assign w_sys_tmp14271 = 32'sh00000070;
	assign w_sys_tmp14273 = (r_run_j_37 - w_sys_tmp14274);
	assign w_sys_tmp14274 = 32'sh0000005f;
	assign w_sys_tmp14276 = (w_sys_tmp14277 + r_run_k_36);
	assign w_sys_tmp14277 = (r_run_copy1_j_361 * w_sys_tmp14278);
	assign w_sys_tmp14278 = 32'sh00000081;
	assign w_sys_tmp14279 = w_sub30_result_dataout;
	assign w_sys_tmp14280 = (w_sys_tmp14281 + r_run_k_36);
	assign w_sys_tmp14281 = (r_run_copy0_j_360 * w_sys_tmp14278);
	assign w_sys_tmp14283 = (r_run_copy0_j_360 + w_sys_intOne);
	assign w_sys_tmp14284 = (r_run_copy1_j_361 + w_sys_intOne);
	assign w_sys_tmp14285 = (r_run_j_37 + w_sys_intOne);
	assign w_sys_tmp14364 = 32'sh00000071;
	assign w_sys_tmp14365 = ( !w_sys_tmp14366 );
	assign w_sys_tmp14366 = (w_sys_tmp14367 < r_run_j_37);
	assign w_sys_tmp14367 = 32'sh00000080;
	assign w_sys_tmp14369 = (r_run_j_37 - w_sys_tmp14370);
	assign w_sys_tmp14370 = 32'sh0000006f;
	assign w_sys_tmp14372 = (w_sys_tmp14373 + r_run_k_36);
	assign w_sys_tmp14373 = (r_run_copy1_j_363 * w_sys_tmp14374);
	assign w_sys_tmp14374 = 32'sh00000081;
	assign w_sys_tmp14375 = w_sub31_result_dataout;
	assign w_sys_tmp14376 = (w_sys_tmp14377 + r_run_k_36);
	assign w_sys_tmp14377 = (r_run_copy0_j_362 * w_sys_tmp14374);
	assign w_sys_tmp14379 = (r_run_copy0_j_362 + w_sys_intOne);
	assign w_sys_tmp14380 = (r_run_copy1_j_363 + w_sys_intOne);
	assign w_sys_tmp14381 = (r_run_j_37 + w_sys_intOne);


	sub19
		sub19_inst(
			.i_fld_T_0_addr_0 (w_sub19_T_addr),
			.i_fld_T_0_datain_0 (w_sub19_T_datain),
			.o_fld_T_0_dataout_0 (w_sub19_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub19_T_r_w),
			.i_fld_U_2_addr_0 (w_sub19_U_addr),
			.i_fld_U_2_datain_0 (w_sub19_U_datain),
			.o_fld_U_2_dataout_0 (w_sub19_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub19_U_r_w),
			.i_fld_V_1_addr_0 (w_sub19_V_addr),
			.i_fld_V_1_datain_0 (w_sub19_V_datain),
			.o_fld_V_1_dataout_0 (w_sub19_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub19_V_r_w),
			.i_fld_result_3_addr_0 (w_sub19_result_addr),
			.i_fld_result_3_datain_0 (w_sub19_result_datain),
			.o_fld_result_3_dataout_0 (w_sub19_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub19_result_r_w),
			.o_run_busy (w_sub19_run_busy),
			.i_run_req (r_sub19_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_T_0_addr_0 (w_sub12_T_addr),
			.i_fld_T_0_datain_0 (w_sub12_T_datain),
			.o_fld_T_0_dataout_0 (w_sub12_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub12_T_r_w),
			.i_fld_U_2_addr_0 (w_sub12_U_addr),
			.i_fld_U_2_datain_0 (w_sub12_U_datain),
			.o_fld_U_2_dataout_0 (w_sub12_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub12_U_r_w),
			.i_fld_V_1_addr_0 (w_sub12_V_addr),
			.i_fld_V_1_datain_0 (w_sub12_V_datain),
			.o_fld_V_1_dataout_0 (w_sub12_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub12_V_r_w),
			.i_fld_result_3_addr_0 (w_sub12_result_addr),
			.i_fld_result_3_datain_0 (w_sub12_result_datain),
			.o_fld_result_3_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub12_result_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_T_0_addr_0 (w_sub11_T_addr),
			.i_fld_T_0_datain_0 (w_sub11_T_datain),
			.o_fld_T_0_dataout_0 (w_sub11_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub11_T_r_w),
			.i_fld_U_2_addr_0 (w_sub11_U_addr),
			.i_fld_U_2_datain_0 (w_sub11_U_datain),
			.o_fld_U_2_dataout_0 (w_sub11_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub11_U_r_w),
			.i_fld_V_1_addr_0 (w_sub11_V_addr),
			.i_fld_V_1_datain_0 (w_sub11_V_datain),
			.o_fld_V_1_dataout_0 (w_sub11_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub11_V_r_w),
			.i_fld_result_3_addr_0 (w_sub11_result_addr),
			.i_fld_result_3_datain_0 (w_sub11_result_datain),
			.o_fld_result_3_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub11_result_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_T_0_addr_0 (w_sub14_T_addr),
			.i_fld_T_0_datain_0 (w_sub14_T_datain),
			.o_fld_T_0_dataout_0 (w_sub14_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub14_T_r_w),
			.i_fld_U_2_addr_0 (w_sub14_U_addr),
			.i_fld_U_2_datain_0 (w_sub14_U_datain),
			.o_fld_U_2_dataout_0 (w_sub14_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub14_U_r_w),
			.i_fld_V_1_addr_0 (w_sub14_V_addr),
			.i_fld_V_1_datain_0 (w_sub14_V_datain),
			.o_fld_V_1_dataout_0 (w_sub14_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub14_V_r_w),
			.i_fld_result_3_addr_0 (w_sub14_result_addr),
			.i_fld_result_3_datain_0 (w_sub14_result_datain),
			.o_fld_result_3_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub14_result_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_T_0_addr_0 (w_sub13_T_addr),
			.i_fld_T_0_datain_0 (w_sub13_T_datain),
			.o_fld_T_0_dataout_0 (w_sub13_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub13_T_r_w),
			.i_fld_U_2_addr_0 (w_sub13_U_addr),
			.i_fld_U_2_datain_0 (w_sub13_U_datain),
			.o_fld_U_2_dataout_0 (w_sub13_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub13_U_r_w),
			.i_fld_V_1_addr_0 (w_sub13_V_addr),
			.i_fld_V_1_datain_0 (w_sub13_V_datain),
			.o_fld_V_1_dataout_0 (w_sub13_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub13_V_r_w),
			.i_fld_result_3_addr_0 (w_sub13_result_addr),
			.i_fld_result_3_datain_0 (w_sub13_result_datain),
			.o_fld_result_3_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub13_result_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub16
		sub16_inst(
			.i_fld_T_0_addr_0 (w_sub16_T_addr),
			.i_fld_T_0_datain_0 (w_sub16_T_datain),
			.o_fld_T_0_dataout_0 (w_sub16_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub16_T_r_w),
			.i_fld_U_2_addr_0 (w_sub16_U_addr),
			.i_fld_U_2_datain_0 (w_sub16_U_datain),
			.o_fld_U_2_dataout_0 (w_sub16_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub16_U_r_w),
			.i_fld_V_1_addr_0 (w_sub16_V_addr),
			.i_fld_V_1_datain_0 (w_sub16_V_datain),
			.o_fld_V_1_dataout_0 (w_sub16_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub16_V_r_w),
			.i_fld_result_3_addr_0 (w_sub16_result_addr),
			.i_fld_result_3_datain_0 (w_sub16_result_datain),
			.o_fld_result_3_dataout_0 (w_sub16_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub16_result_r_w),
			.o_run_busy (w_sub16_run_busy),
			.i_run_req (r_sub16_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_T_0_addr_0 (w_sub15_T_addr),
			.i_fld_T_0_datain_0 (w_sub15_T_datain),
			.o_fld_T_0_dataout_0 (w_sub15_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub15_T_r_w),
			.i_fld_U_2_addr_0 (w_sub15_U_addr),
			.i_fld_U_2_datain_0 (w_sub15_U_datain),
			.o_fld_U_2_dataout_0 (w_sub15_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub15_U_r_w),
			.i_fld_V_1_addr_0 (w_sub15_V_addr),
			.i_fld_V_1_datain_0 (w_sub15_V_datain),
			.o_fld_V_1_dataout_0 (w_sub15_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub15_V_r_w),
			.i_fld_result_3_addr_0 (w_sub15_result_addr),
			.i_fld_result_3_datain_0 (w_sub15_result_datain),
			.o_fld_result_3_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub15_result_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub18
		sub18_inst(
			.i_fld_T_0_addr_0 (w_sub18_T_addr),
			.i_fld_T_0_datain_0 (w_sub18_T_datain),
			.o_fld_T_0_dataout_0 (w_sub18_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub18_T_r_w),
			.i_fld_U_2_addr_0 (w_sub18_U_addr),
			.i_fld_U_2_datain_0 (w_sub18_U_datain),
			.o_fld_U_2_dataout_0 (w_sub18_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub18_U_r_w),
			.i_fld_V_1_addr_0 (w_sub18_V_addr),
			.i_fld_V_1_datain_0 (w_sub18_V_datain),
			.o_fld_V_1_dataout_0 (w_sub18_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub18_V_r_w),
			.i_fld_result_3_addr_0 (w_sub18_result_addr),
			.i_fld_result_3_datain_0 (w_sub18_result_datain),
			.o_fld_result_3_dataout_0 (w_sub18_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub18_result_r_w),
			.o_run_busy (w_sub18_run_busy),
			.i_run_req (r_sub18_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub17
		sub17_inst(
			.i_fld_T_0_addr_0 (w_sub17_T_addr),
			.i_fld_T_0_datain_0 (w_sub17_T_datain),
			.o_fld_T_0_dataout_0 (w_sub17_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub17_T_r_w),
			.i_fld_U_2_addr_0 (w_sub17_U_addr),
			.i_fld_U_2_datain_0 (w_sub17_U_datain),
			.o_fld_U_2_dataout_0 (w_sub17_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub17_U_r_w),
			.i_fld_V_1_addr_0 (w_sub17_V_addr),
			.i_fld_V_1_datain_0 (w_sub17_V_datain),
			.o_fld_V_1_dataout_0 (w_sub17_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub17_V_r_w),
			.i_fld_result_3_addr_0 (w_sub17_result_addr),
			.i_fld_result_3_datain_0 (w_sub17_result_datain),
			.o_fld_result_3_dataout_0 (w_sub17_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub17_result_r_w),
			.o_run_busy (w_sub17_run_busy),
			.i_run_req (r_sub17_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub20
		sub20_inst(
			.i_fld_T_0_addr_0 (w_sub20_T_addr),
			.i_fld_T_0_datain_0 (w_sub20_T_datain),
			.o_fld_T_0_dataout_0 (w_sub20_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub20_T_r_w),
			.i_fld_U_2_addr_0 (w_sub20_U_addr),
			.i_fld_U_2_datain_0 (w_sub20_U_datain),
			.o_fld_U_2_dataout_0 (w_sub20_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub20_U_r_w),
			.i_fld_V_1_addr_0 (w_sub20_V_addr),
			.i_fld_V_1_datain_0 (w_sub20_V_datain),
			.o_fld_V_1_dataout_0 (w_sub20_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub20_V_r_w),
			.i_fld_result_3_addr_0 (w_sub20_result_addr),
			.i_fld_result_3_datain_0 (w_sub20_result_datain),
			.o_fld_result_3_dataout_0 (w_sub20_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub20_result_r_w),
			.o_run_busy (w_sub20_run_busy),
			.i_run_req (r_sub20_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub21
		sub21_inst(
			.i_fld_T_0_addr_0 (w_sub21_T_addr),
			.i_fld_T_0_datain_0 (w_sub21_T_datain),
			.o_fld_T_0_dataout_0 (w_sub21_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub21_T_r_w),
			.i_fld_U_2_addr_0 (w_sub21_U_addr),
			.i_fld_U_2_datain_0 (w_sub21_U_datain),
			.o_fld_U_2_dataout_0 (w_sub21_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub21_U_r_w),
			.i_fld_V_1_addr_0 (w_sub21_V_addr),
			.i_fld_V_1_datain_0 (w_sub21_V_datain),
			.o_fld_V_1_dataout_0 (w_sub21_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub21_V_r_w),
			.i_fld_result_3_addr_0 (w_sub21_result_addr),
			.i_fld_result_3_datain_0 (w_sub21_result_datain),
			.o_fld_result_3_dataout_0 (w_sub21_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub21_result_r_w),
			.o_run_busy (w_sub21_run_busy),
			.i_run_req (r_sub21_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub28
		sub28_inst(
			.i_fld_T_0_addr_0 (w_sub28_T_addr),
			.i_fld_T_0_datain_0 (w_sub28_T_datain),
			.o_fld_T_0_dataout_0 (w_sub28_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub28_T_r_w),
			.i_fld_U_2_addr_0 (w_sub28_U_addr),
			.i_fld_U_2_datain_0 (w_sub28_U_datain),
			.o_fld_U_2_dataout_0 (w_sub28_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub28_U_r_w),
			.i_fld_V_1_addr_0 (w_sub28_V_addr),
			.i_fld_V_1_datain_0 (w_sub28_V_datain),
			.o_fld_V_1_dataout_0 (w_sub28_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub28_V_r_w),
			.i_fld_result_3_addr_0 (w_sub28_result_addr),
			.i_fld_result_3_datain_0 (w_sub28_result_datain),
			.o_fld_result_3_dataout_0 (w_sub28_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub28_result_r_w),
			.o_run_busy (w_sub28_run_busy),
			.i_run_req (r_sub28_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub29
		sub29_inst(
			.i_fld_T_0_addr_0 (w_sub29_T_addr),
			.i_fld_T_0_datain_0 (w_sub29_T_datain),
			.o_fld_T_0_dataout_0 (w_sub29_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub29_T_r_w),
			.i_fld_U_2_addr_0 (w_sub29_U_addr),
			.i_fld_U_2_datain_0 (w_sub29_U_datain),
			.o_fld_U_2_dataout_0 (w_sub29_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub29_U_r_w),
			.i_fld_V_1_addr_0 (w_sub29_V_addr),
			.i_fld_V_1_datain_0 (w_sub29_V_datain),
			.o_fld_V_1_dataout_0 (w_sub29_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub29_V_r_w),
			.i_fld_result_3_addr_0 (w_sub29_result_addr),
			.i_fld_result_3_datain_0 (w_sub29_result_datain),
			.o_fld_result_3_dataout_0 (w_sub29_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub29_result_r_w),
			.o_run_busy (w_sub29_run_busy),
			.i_run_req (r_sub29_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub26
		sub26_inst(
			.i_fld_T_0_addr_0 (w_sub26_T_addr),
			.i_fld_T_0_datain_0 (w_sub26_T_datain),
			.o_fld_T_0_dataout_0 (w_sub26_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub26_T_r_w),
			.i_fld_U_2_addr_0 (w_sub26_U_addr),
			.i_fld_U_2_datain_0 (w_sub26_U_datain),
			.o_fld_U_2_dataout_0 (w_sub26_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub26_U_r_w),
			.i_fld_V_1_addr_0 (w_sub26_V_addr),
			.i_fld_V_1_datain_0 (w_sub26_V_datain),
			.o_fld_V_1_dataout_0 (w_sub26_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub26_V_r_w),
			.i_fld_result_3_addr_0 (w_sub26_result_addr),
			.i_fld_result_3_datain_0 (w_sub26_result_datain),
			.o_fld_result_3_dataout_0 (w_sub26_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub26_result_r_w),
			.o_run_busy (w_sub26_run_busy),
			.i_run_req (r_sub26_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub09
		sub09_inst(
			.i_fld_T_0_addr_0 (w_sub09_T_addr),
			.i_fld_T_0_datain_0 (w_sub09_T_datain),
			.o_fld_T_0_dataout_0 (w_sub09_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub09_T_r_w),
			.i_fld_U_2_addr_0 (w_sub09_U_addr),
			.i_fld_U_2_datain_0 (w_sub09_U_datain),
			.o_fld_U_2_dataout_0 (w_sub09_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub09_U_r_w),
			.i_fld_V_1_addr_0 (w_sub09_V_addr),
			.i_fld_V_1_datain_0 (w_sub09_V_datain),
			.o_fld_V_1_dataout_0 (w_sub09_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub09_V_r_w),
			.i_fld_result_3_addr_0 (w_sub09_result_addr),
			.i_fld_result_3_datain_0 (w_sub09_result_datain),
			.o_fld_result_3_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub09_result_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub27
		sub27_inst(
			.i_fld_T_0_addr_0 (w_sub27_T_addr),
			.i_fld_T_0_datain_0 (w_sub27_T_datain),
			.o_fld_T_0_dataout_0 (w_sub27_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub27_T_r_w),
			.i_fld_U_2_addr_0 (w_sub27_U_addr),
			.i_fld_U_2_datain_0 (w_sub27_U_datain),
			.o_fld_U_2_dataout_0 (w_sub27_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub27_U_r_w),
			.i_fld_V_1_addr_0 (w_sub27_V_addr),
			.i_fld_V_1_datain_0 (w_sub27_V_datain),
			.o_fld_V_1_dataout_0 (w_sub27_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub27_V_r_w),
			.i_fld_result_3_addr_0 (w_sub27_result_addr),
			.i_fld_result_3_datain_0 (w_sub27_result_datain),
			.o_fld_result_3_dataout_0 (w_sub27_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub27_result_r_w),
			.o_run_busy (w_sub27_run_busy),
			.i_run_req (r_sub27_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_T_0_addr_0 (w_sub08_T_addr),
			.i_fld_T_0_datain_0 (w_sub08_T_datain),
			.o_fld_T_0_dataout_0 (w_sub08_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub08_T_r_w),
			.i_fld_U_2_addr_0 (w_sub08_U_addr),
			.i_fld_U_2_datain_0 (w_sub08_U_datain),
			.o_fld_U_2_dataout_0 (w_sub08_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub08_U_r_w),
			.i_fld_V_1_addr_0 (w_sub08_V_addr),
			.i_fld_V_1_datain_0 (w_sub08_V_datain),
			.o_fld_V_1_dataout_0 (w_sub08_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub08_V_r_w),
			.i_fld_result_3_addr_0 (w_sub08_result_addr),
			.i_fld_result_3_datain_0 (w_sub08_result_datain),
			.o_fld_result_3_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub08_result_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub24
		sub24_inst(
			.i_fld_T_0_addr_0 (w_sub24_T_addr),
			.i_fld_T_0_datain_0 (w_sub24_T_datain),
			.o_fld_T_0_dataout_0 (w_sub24_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub24_T_r_w),
			.i_fld_U_2_addr_0 (w_sub24_U_addr),
			.i_fld_U_2_datain_0 (w_sub24_U_datain),
			.o_fld_U_2_dataout_0 (w_sub24_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub24_U_r_w),
			.i_fld_V_1_addr_0 (w_sub24_V_addr),
			.i_fld_V_1_datain_0 (w_sub24_V_datain),
			.o_fld_V_1_dataout_0 (w_sub24_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub24_V_r_w),
			.i_fld_result_3_addr_0 (w_sub24_result_addr),
			.i_fld_result_3_datain_0 (w_sub24_result_datain),
			.o_fld_result_3_dataout_0 (w_sub24_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub24_result_r_w),
			.o_run_busy (w_sub24_run_busy),
			.i_run_req (r_sub24_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub25
		sub25_inst(
			.i_fld_T_0_addr_0 (w_sub25_T_addr),
			.i_fld_T_0_datain_0 (w_sub25_T_datain),
			.o_fld_T_0_dataout_0 (w_sub25_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub25_T_r_w),
			.i_fld_U_2_addr_0 (w_sub25_U_addr),
			.i_fld_U_2_datain_0 (w_sub25_U_datain),
			.o_fld_U_2_dataout_0 (w_sub25_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub25_U_r_w),
			.i_fld_V_1_addr_0 (w_sub25_V_addr),
			.i_fld_V_1_datain_0 (w_sub25_V_datain),
			.o_fld_V_1_dataout_0 (w_sub25_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub25_V_r_w),
			.i_fld_result_3_addr_0 (w_sub25_result_addr),
			.i_fld_result_3_datain_0 (w_sub25_result_datain),
			.o_fld_result_3_dataout_0 (w_sub25_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub25_result_r_w),
			.o_run_busy (w_sub25_run_busy),
			.i_run_req (r_sub25_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub22
		sub22_inst(
			.i_fld_T_0_addr_0 (w_sub22_T_addr),
			.i_fld_T_0_datain_0 (w_sub22_T_datain),
			.o_fld_T_0_dataout_0 (w_sub22_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub22_T_r_w),
			.i_fld_U_2_addr_0 (w_sub22_U_addr),
			.i_fld_U_2_datain_0 (w_sub22_U_datain),
			.o_fld_U_2_dataout_0 (w_sub22_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub22_U_r_w),
			.i_fld_V_1_addr_0 (w_sub22_V_addr),
			.i_fld_V_1_datain_0 (w_sub22_V_datain),
			.o_fld_V_1_dataout_0 (w_sub22_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub22_V_r_w),
			.i_fld_result_3_addr_0 (w_sub22_result_addr),
			.i_fld_result_3_datain_0 (w_sub22_result_datain),
			.o_fld_result_3_dataout_0 (w_sub22_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub22_result_r_w),
			.o_run_busy (w_sub22_run_busy),
			.i_run_req (r_sub22_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub23
		sub23_inst(
			.i_fld_T_0_addr_0 (w_sub23_T_addr),
			.i_fld_T_0_datain_0 (w_sub23_T_datain),
			.o_fld_T_0_dataout_0 (w_sub23_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub23_T_r_w),
			.i_fld_U_2_addr_0 (w_sub23_U_addr),
			.i_fld_U_2_datain_0 (w_sub23_U_datain),
			.o_fld_U_2_dataout_0 (w_sub23_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub23_U_r_w),
			.i_fld_V_1_addr_0 (w_sub23_V_addr),
			.i_fld_V_1_datain_0 (w_sub23_V_datain),
			.o_fld_V_1_dataout_0 (w_sub23_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub23_V_r_w),
			.i_fld_result_3_addr_0 (w_sub23_result_addr),
			.i_fld_result_3_datain_0 (w_sub23_result_datain),
			.o_fld_result_3_dataout_0 (w_sub23_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub23_result_r_w),
			.o_run_busy (w_sub23_run_busy),
			.i_run_req (r_sub23_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_T_0_addr_0 (w_sub03_T_addr),
			.i_fld_T_0_datain_0 (w_sub03_T_datain),
			.o_fld_T_0_dataout_0 (w_sub03_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub03_T_r_w),
			.i_fld_U_2_addr_0 (w_sub03_U_addr),
			.i_fld_U_2_datain_0 (w_sub03_U_datain),
			.o_fld_U_2_dataout_0 (w_sub03_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub03_U_r_w),
			.i_fld_V_1_addr_0 (w_sub03_V_addr),
			.i_fld_V_1_datain_0 (w_sub03_V_datain),
			.o_fld_V_1_dataout_0 (w_sub03_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub03_V_r_w),
			.i_fld_result_3_addr_0 (w_sub03_result_addr),
			.i_fld_result_3_datain_0 (w_sub03_result_datain),
			.o_fld_result_3_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub03_result_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_T_0_addr_0 (w_sub02_T_addr),
			.i_fld_T_0_datain_0 (w_sub02_T_datain),
			.o_fld_T_0_dataout_0 (w_sub02_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub02_T_r_w),
			.i_fld_U_2_addr_0 (w_sub02_U_addr),
			.i_fld_U_2_datain_0 (w_sub02_U_datain),
			.o_fld_U_2_dataout_0 (w_sub02_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub02_U_r_w),
			.i_fld_V_1_addr_0 (w_sub02_V_addr),
			.i_fld_V_1_datain_0 (w_sub02_V_datain),
			.o_fld_V_1_dataout_0 (w_sub02_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub02_V_r_w),
			.i_fld_result_3_addr_0 (w_sub02_result_addr),
			.i_fld_result_3_datain_0 (w_sub02_result_datain),
			.o_fld_result_3_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub02_result_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_T_0_addr_0 (w_sub01_T_addr),
			.i_fld_T_0_datain_0 (w_sub01_T_datain),
			.o_fld_T_0_dataout_0 (w_sub01_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub01_T_r_w),
			.i_fld_U_2_addr_0 (w_sub01_U_addr),
			.i_fld_U_2_datain_0 (w_sub01_U_datain),
			.o_fld_U_2_dataout_0 (w_sub01_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub01_U_r_w),
			.i_fld_V_1_addr_0 (w_sub01_V_addr),
			.i_fld_V_1_datain_0 (w_sub01_V_datain),
			.o_fld_V_1_dataout_0 (w_sub01_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub01_V_r_w),
			.i_fld_result_3_addr_0 (w_sub01_result_addr),
			.i_fld_result_3_datain_0 (w_sub01_result_datain),
			.o_fld_result_3_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub01_result_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_T_0_addr_0 (w_sub00_T_addr),
			.i_fld_T_0_datain_0 (w_sub00_T_datain),
			.o_fld_T_0_dataout_0 (w_sub00_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub00_T_r_w),
			.i_fld_U_2_addr_0 (w_sub00_U_addr),
			.i_fld_U_2_datain_0 (w_sub00_U_datain),
			.o_fld_U_2_dataout_0 (w_sub00_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub00_U_r_w),
			.i_fld_V_1_addr_0 (w_sub00_V_addr),
			.i_fld_V_1_datain_0 (w_sub00_V_datain),
			.o_fld_V_1_dataout_0 (w_sub00_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub00_V_r_w),
			.i_fld_result_3_addr_0 (w_sub00_result_addr),
			.i_fld_result_3_datain_0 (w_sub00_result_datain),
			.o_fld_result_3_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub00_result_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_T_0_addr_0 (w_sub07_T_addr),
			.i_fld_T_0_datain_0 (w_sub07_T_datain),
			.o_fld_T_0_dataout_0 (w_sub07_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub07_T_r_w),
			.i_fld_U_2_addr_0 (w_sub07_U_addr),
			.i_fld_U_2_datain_0 (w_sub07_U_datain),
			.o_fld_U_2_dataout_0 (w_sub07_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub07_U_r_w),
			.i_fld_V_1_addr_0 (w_sub07_V_addr),
			.i_fld_V_1_datain_0 (w_sub07_V_datain),
			.o_fld_V_1_dataout_0 (w_sub07_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub07_V_r_w),
			.i_fld_result_3_addr_0 (w_sub07_result_addr),
			.i_fld_result_3_datain_0 (w_sub07_result_datain),
			.o_fld_result_3_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub07_result_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_T_0_addr_0 (w_sub06_T_addr),
			.i_fld_T_0_datain_0 (w_sub06_T_datain),
			.o_fld_T_0_dataout_0 (w_sub06_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub06_T_r_w),
			.i_fld_U_2_addr_0 (w_sub06_U_addr),
			.i_fld_U_2_datain_0 (w_sub06_U_datain),
			.o_fld_U_2_dataout_0 (w_sub06_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub06_U_r_w),
			.i_fld_V_1_addr_0 (w_sub06_V_addr),
			.i_fld_V_1_datain_0 (w_sub06_V_datain),
			.o_fld_V_1_dataout_0 (w_sub06_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub06_V_r_w),
			.i_fld_result_3_addr_0 (w_sub06_result_addr),
			.i_fld_result_3_datain_0 (w_sub06_result_datain),
			.o_fld_result_3_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub06_result_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_T_0_addr_0 (w_sub05_T_addr),
			.i_fld_T_0_datain_0 (w_sub05_T_datain),
			.o_fld_T_0_dataout_0 (w_sub05_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub05_T_r_w),
			.i_fld_U_2_addr_0 (w_sub05_U_addr),
			.i_fld_U_2_datain_0 (w_sub05_U_datain),
			.o_fld_U_2_dataout_0 (w_sub05_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub05_U_r_w),
			.i_fld_V_1_addr_0 (w_sub05_V_addr),
			.i_fld_V_1_datain_0 (w_sub05_V_datain),
			.o_fld_V_1_dataout_0 (w_sub05_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub05_V_r_w),
			.i_fld_result_3_addr_0 (w_sub05_result_addr),
			.i_fld_result_3_datain_0 (w_sub05_result_datain),
			.o_fld_result_3_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub05_result_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_T_0_addr_0 (w_sub04_T_addr),
			.i_fld_T_0_datain_0 (w_sub04_T_datain),
			.o_fld_T_0_dataout_0 (w_sub04_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub04_T_r_w),
			.i_fld_U_2_addr_0 (w_sub04_U_addr),
			.i_fld_U_2_datain_0 (w_sub04_U_datain),
			.o_fld_U_2_dataout_0 (w_sub04_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub04_U_r_w),
			.i_fld_V_1_addr_0 (w_sub04_V_addr),
			.i_fld_V_1_datain_0 (w_sub04_V_datain),
			.o_fld_V_1_dataout_0 (w_sub04_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub04_V_r_w),
			.i_fld_result_3_addr_0 (w_sub04_result_addr),
			.i_fld_result_3_datain_0 (w_sub04_result_datain),
			.o_fld_result_3_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub04_result_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_T_0_addr_0 (w_sub10_T_addr),
			.i_fld_T_0_datain_0 (w_sub10_T_datain),
			.o_fld_T_0_dataout_0 (w_sub10_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub10_T_r_w),
			.i_fld_U_2_addr_0 (w_sub10_U_addr),
			.i_fld_U_2_datain_0 (w_sub10_U_datain),
			.o_fld_U_2_dataout_0 (w_sub10_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub10_U_r_w),
			.i_fld_V_1_addr_0 (w_sub10_V_addr),
			.i_fld_V_1_datain_0 (w_sub10_V_datain),
			.o_fld_V_1_dataout_0 (w_sub10_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub10_V_r_w),
			.i_fld_result_3_addr_0 (w_sub10_result_addr),
			.i_fld_result_3_datain_0 (w_sub10_result_datain),
			.o_fld_result_3_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub10_result_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub31
		sub31_inst(
			.i_fld_T_0_addr_0 (w_sub31_T_addr),
			.i_fld_T_0_datain_0 (w_sub31_T_datain),
			.o_fld_T_0_dataout_0 (w_sub31_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub31_T_r_w),
			.i_fld_U_2_addr_0 (w_sub31_U_addr),
			.i_fld_U_2_datain_0 (w_sub31_U_datain),
			.o_fld_U_2_dataout_0 (w_sub31_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub31_U_r_w),
			.i_fld_V_1_addr_0 (w_sub31_V_addr),
			.i_fld_V_1_datain_0 (w_sub31_V_datain),
			.o_fld_V_1_dataout_0 (w_sub31_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub31_V_r_w),
			.i_fld_result_3_addr_0 (w_sub31_result_addr),
			.i_fld_result_3_datain_0 (w_sub31_result_datain),
			.o_fld_result_3_dataout_0 (w_sub31_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub31_result_r_w),
			.o_run_busy (w_sub31_run_busy),
			.i_run_req (r_sub31_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub30
		sub30_inst(
			.i_fld_T_0_addr_0 (w_sub30_T_addr),
			.i_fld_T_0_datain_0 (w_sub30_T_datain),
			.o_fld_T_0_dataout_0 (w_sub30_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub30_T_r_w),
			.i_fld_U_2_addr_0 (w_sub30_U_addr),
			.i_fld_U_2_datain_0 (w_sub30_U_datain),
			.o_fld_U_2_dataout_0 (w_sub30_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub30_U_r_w),
			.i_fld_V_1_addr_0 (w_sub30_V_addr),
			.i_fld_V_1_datain_0 (w_sub30_V_datain),
			.o_fld_V_1_dataout_0 (w_sub30_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub30_V_r_w),
			.i_fld_result_3_addr_0 (w_sub30_result_addr),
			.i_fld_result_3_datain_0 (w_sub30_result_datain),
			.o_fld_result_3_dataout_0 (w_sub30_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub30_result_r_w),
			.o_run_busy (w_sub30_run_busy),
			.i_run_req (r_sub30_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_V_3(
			.clk (clock),
			.ce_0 (w_fld_V_3_ce_0),
			.addr_0 (w_fld_V_3_addr_0),
			.datain_0 (w_fld_V_3_datain_0),
			.dataout_0 (w_fld_V_3_dataout_0),
			.r_w_0 (w_fld_V_3_r_w_0),
			.ce_1 (w_fld_V_3_ce_1),
			.addr_1 (r_fld_V_3_addr_1),
			.datain_1 (r_fld_V_3_datain_1),
			.dataout_1 (w_fld_V_3_dataout_1),
			.r_w_1 (r_fld_V_3_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp38;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==6'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1b)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp18;

									end
									else
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
									else
									if((6'h7<=r_sys_run_step && r_sys_run_step<=6'hb) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'hf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_43;

									end
									else
									if((r_sys_run_step==6'h18)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h16)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp36;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp37;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h16)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_48;

									end
									else
									if((6'h7<=r_sys_run_step && r_sys_run_step<=6'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h13) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						10'h207: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 10'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h0: begin
							r_sys_run_phase <= 10'h2;
						end

						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h4;

									end
								end

							endcase
						end

						10'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h5;

									end
								end

							endcase
						end

						10'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12) ? 10'h9 : 10'hf);

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h5;

									end
								end

							endcase
						end

						10'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'ha;

									end
								end

							endcase
						end

						10'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp15) ? 10'hd : 10'h6);

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_phase <= 10'ha;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h10;

									end
								end

							endcase
						end

						10'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp226) ? 10'h14 : 10'h44);

									end
								end

							endcase
						end

						10'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h10;

									end
								end

							endcase
						end

						10'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h15;

									end
								end

							endcase
						end

						10'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp230) ? 10'h18 : 10'h1a);

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h15;

									end
								end

							endcase
						end

						10'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1b;

									end
								end

							endcase
						end

						10'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp445) ? 10'h1e : 10'h20);

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1b;

									end
								end

							endcase
						end

						10'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h21;

									end
								end

							endcase
						end

						10'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp660) ? 10'h24 : 10'h26);

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h21;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h27;

									end
								end

							endcase
						end

						10'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp875) ? 10'h2a : 10'h2c);

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h27;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h2d;

									end
								end

							endcase
						end

						10'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1090) ? 10'h30 : 10'h32);

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h2d;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h33;

									end
								end

							endcase
						end

						10'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1305) ? 10'h36 : 10'h38);

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h33;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h39;

									end
								end

							endcase
						end

						10'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1520) ? 10'h3c : 10'h3e);

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h39;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h3f;

									end
								end

							endcase
						end

						10'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1735) ? 10'h42 : 10'h11);

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h3f;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h45;

									end
								end

							endcase
						end

						10'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1949) ? 10'h49 : 10'h79);

									end
								end

							endcase
						end

						10'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h45;

									end
								end

							endcase
						end

						10'h49: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h4a;

									end
								end

							endcase
						end

						10'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1953) ? 10'h4d : 10'h4f);

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h4a;

									end
								end

							endcase
						end

						10'h4f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h50;

									end
								end

							endcase
						end

						10'h50: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2168) ? 10'h53 : 10'h55);

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h50;

									end
								end

							endcase
						end

						10'h55: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h56;

									end
								end

							endcase
						end

						10'h56: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2383) ? 10'h59 : 10'h5b);

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h56;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h5c;

									end
								end

							endcase
						end

						10'h5c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2598) ? 10'h5f : 10'h61);

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h5c;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h62;

									end
								end

							endcase
						end

						10'h62: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2813) ? 10'h65 : 10'h67);

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h62;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h68;

									end
								end

							endcase
						end

						10'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3028) ? 10'h6b : 10'h6d);

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h68;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h6e;

									end
								end

							endcase
						end

						10'h6e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3243) ? 10'h71 : 10'h73);

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h6e;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h74;

									end
								end

							endcase
						end

						10'h74: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3458) ? 10'h77 : 10'h46);

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h74;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h7a;

									end
								end

							endcase
						end

						10'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3672) ? 10'h7e : 10'hae);

									end
								end

							endcase
						end

						10'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h7a;

									end
								end

							endcase
						end

						10'h7e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h7f;

									end
								end

							endcase
						end

						10'h7f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3676) ? 10'h82 : 10'h84);

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h7f;

									end
								end

							endcase
						end

						10'h84: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h85;

									end
								end

							endcase
						end

						10'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3891) ? 10'h88 : 10'h8a);

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h85;

									end
								end

							endcase
						end

						10'h8a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h8b;

									end
								end

							endcase
						end

						10'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4106) ? 10'h8e : 10'h90);

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h8b;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h91;

									end
								end

							endcase
						end

						10'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4321) ? 10'h94 : 10'h96);

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h91;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h97;

									end
								end

							endcase
						end

						10'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4536) ? 10'h9a : 10'h9c);

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h97;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h9d;

									end
								end

							endcase
						end

						10'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4751) ? 10'ha0 : 10'ha2);

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h9d;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'ha3;

									end
								end

							endcase
						end

						10'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4966) ? 10'ha6 : 10'ha8);

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'ha3;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'ha9;

									end
								end

							endcase
						end

						10'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5181) ? 10'hac : 10'h7b);

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'ha9;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'haf;

									end
								end

							endcase
						end

						10'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5395) ? 10'hb3 : 10'he3);

									end
								end

							endcase
						end

						10'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'haf;

									end
								end

							endcase
						end

						10'hb3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hb4;

									end
								end

							endcase
						end

						10'hb4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5399) ? 10'hb7 : 10'hb9);

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hb4;

									end
								end

							endcase
						end

						10'hb9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hba;

									end
								end

							endcase
						end

						10'hba: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5614) ? 10'hbd : 10'hbf);

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hba;

									end
								end

							endcase
						end

						10'hbf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hc0;

									end
								end

							endcase
						end

						10'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5829) ? 10'hc3 : 10'hc5);

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hc0;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hc6;

									end
								end

							endcase
						end

						10'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6044) ? 10'hc9 : 10'hcb);

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hc6;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hcc;

									end
								end

							endcase
						end

						10'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6259) ? 10'hcf : 10'hd1);

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hcc;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hd2;

									end
								end

							endcase
						end

						10'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6474) ? 10'hd5 : 10'hd7);

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hd2;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hd8;

									end
								end

							endcase
						end

						10'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6689) ? 10'hdb : 10'hdd);

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hd8;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hde;

									end
								end

							endcase
						end

						10'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6904) ? 10'he1 : 10'hb0);

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hde;

									end
								end

							endcase
						end

						10'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'he4;

									end
								end

							endcase
						end

						10'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7118) ? 10'he7 : 10'h133);

									end
								end

							endcase
						end

						10'he5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'he4;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 10'he9;

									end
								end

							endcase
						end

						10'he9: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 10'heb;

									end
								end

							endcase
						end

						10'heb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hec;

									end
								end

							endcase
						end

						10'hec: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7122) ? 10'hef : 10'hf1);

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'hec;

									end
								end

							endcase
						end

						10'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hf2;

									end
								end

							endcase
						end

						10'hf2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7206) ? 10'hf5 : 10'hf7);

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'hf2;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hf8;

									end
								end

							endcase
						end

						10'hf8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7290) ? 10'hfb : 10'hfd);

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'hf8;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hfe;

									end
								end

							endcase
						end

						10'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7374) ? 10'h101 : 10'h103);

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'hfe;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h104;

									end
								end

							endcase
						end

						10'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7457) ? 10'h107 : 10'h109);

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h104;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h10a;

									end
								end

							endcase
						end

						10'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7958) ? 10'h10d : 10'h10f);

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h10a;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h110;

									end
								end

							endcase
						end

						10'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8459) ? 10'h113 : 10'h115);

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h110;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h116;

									end
								end

							endcase
						end

						10'h116: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8960) ? 10'h119 : 10'h11b);

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h116;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h11c;

									end
								end

							endcase
						end

						10'h11c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9461) ? 10'h11f : 10'h121);

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h11c;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h122;

									end
								end

							endcase
						end

						10'h122: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9962) ? 10'h125 : 10'h127);

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h122;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h128;

									end
								end

							endcase
						end

						10'h128: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10463) ? 10'h12b : 10'h12d);

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h128;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h12e;

									end
								end

							endcase
						end

						10'h12e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10964) ? 10'h131 : 10'he5);

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3a)) begin
										r_sys_run_phase <= 10'h12e;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h134;

									end
								end

							endcase
						end

						10'h134: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11453) ? 10'h138 : 10'h168);

									end
								end

							endcase
						end

						10'h135: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h134;

									end
								end

							endcase
						end

						10'h138: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h139;

									end
								end

							endcase
						end

						10'h139: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11458) ? 10'h13c : 10'h13e);

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h139;

									end
								end

							endcase
						end

						10'h13e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h13f;

									end
								end

							endcase
						end

						10'h13f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11533) ? 10'h142 : 10'h144);

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h13f;

									end
								end

							endcase
						end

						10'h144: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h145;

									end
								end

							endcase
						end

						10'h145: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11629) ? 10'h148 : 10'h14a);

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h145;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h14b;

									end
								end

							endcase
						end

						10'h14b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11725) ? 10'h14e : 10'h150);

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h14b;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h151;

									end
								end

							endcase
						end

						10'h151: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11821) ? 10'h154 : 10'h156);

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h151;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h157;

									end
								end

							endcase
						end

						10'h157: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp11917) ? 10'h15a : 10'h15c);

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h157;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h15d;

									end
								end

							endcase
						end

						10'h15d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12013) ? 10'h160 : 10'h162);

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h15d;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h163;

									end
								end

							endcase
						end

						10'h163: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12109) ? 10'h166 : 10'h135);

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h163;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h169;

									end
								end

							endcase
						end

						10'h169: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12205) ? 10'h16d : 10'h19d);

									end
								end

							endcase
						end

						10'h16a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h169;

									end
								end

							endcase
						end

						10'h16d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h16e;

									end
								end

							endcase
						end

						10'h16e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12210) ? 10'h171 : 10'h173);

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h16e;

									end
								end

							endcase
						end

						10'h173: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h174;

									end
								end

							endcase
						end

						10'h174: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12285) ? 10'h177 : 10'h179);

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h174;

									end
								end

							endcase
						end

						10'h179: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h17a;

									end
								end

							endcase
						end

						10'h17a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12381) ? 10'h17d : 10'h17f);

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h17a;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h180;

									end
								end

							endcase
						end

						10'h180: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12477) ? 10'h183 : 10'h185);

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h180;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h186;

									end
								end

							endcase
						end

						10'h186: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12573) ? 10'h189 : 10'h18b);

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h186;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h18c;

									end
								end

							endcase
						end

						10'h18c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12669) ? 10'h18f : 10'h191);

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h18c;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h192;

									end
								end

							endcase
						end

						10'h192: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12765) ? 10'h195 : 10'h197);

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h192;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h198;

									end
								end

							endcase
						end

						10'h198: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12861) ? 10'h19b : 10'h16a);

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h198;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h19e;

									end
								end

							endcase
						end

						10'h19e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12957) ? 10'h1a2 : 10'h1d2);

									end
								end

							endcase
						end

						10'h19f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h19e;

									end
								end

							endcase
						end

						10'h1a2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1a3;

									end
								end

							endcase
						end

						10'h1a3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12962) ? 10'h1a6 : 10'h1a8);

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1a3;

									end
								end

							endcase
						end

						10'h1a8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1a9;

									end
								end

							endcase
						end

						10'h1a9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13037) ? 10'h1ac : 10'h1ae);

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1a9;

									end
								end

							endcase
						end

						10'h1ae: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1af;

									end
								end

							endcase
						end

						10'h1af: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13133) ? 10'h1b2 : 10'h1b4);

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1af;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1b5;

									end
								end

							endcase
						end

						10'h1b5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13229) ? 10'h1b8 : 10'h1ba);

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1b5;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1bb;

									end
								end

							endcase
						end

						10'h1bb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13325) ? 10'h1be : 10'h1c0);

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1bb;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1c1;

									end
								end

							endcase
						end

						10'h1c1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13421) ? 10'h1c4 : 10'h1c6);

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1c1;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1c7;

									end
								end

							endcase
						end

						10'h1c7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13517) ? 10'h1ca : 10'h1cc);

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1c7;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1cd;

									end
								end

							endcase
						end

						10'h1cd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13613) ? 10'h1d0 : 10'h19f);

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1cd;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1d3;

									end
								end

							endcase
						end

						10'h1d3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13709) ? 10'h1d7 : 10'h207);

									end
								end

							endcase
						end

						10'h1d4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1d3;

									end
								end

							endcase
						end

						10'h1d7: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1d8;

									end
								end

							endcase
						end

						10'h1d8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13714) ? 10'h1db : 10'h1dd);

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1d8;

									end
								end

							endcase
						end

						10'h1dd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1de;

									end
								end

							endcase
						end

						10'h1de: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13789) ? 10'h1e1 : 10'h1e3);

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1de;

									end
								end

							endcase
						end

						10'h1e3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1e4;

									end
								end

							endcase
						end

						10'h1e4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13885) ? 10'h1e7 : 10'h1e9);

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1e4;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1ea;

									end
								end

							endcase
						end

						10'h1ea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13981) ? 10'h1ed : 10'h1ef);

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1ea;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1f0;

									end
								end

							endcase
						end

						10'h1f0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp14077) ? 10'h1f3 : 10'h1f5);

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1f0;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1f6;

									end
								end

							endcase
						end

						10'h1f6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp14173) ? 10'h1f9 : 10'h1fb);

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1f6;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1fc;

									end
								end

							endcase
						end

						10'h1fc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp14269) ? 10'h1ff : 10'h201);

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1fc;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h202;

									end
								end

							endcase
						end

						10'h202: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp14365) ? 10'h205 : 10'h1d4);

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h202;

									end
								end

							endcase
						end

						10'h207: begin
							r_sys_run_phase <= 10'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h50: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h56: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h5c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h62: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h6e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h74: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h7f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h8a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hb4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hba: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hbf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'he5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'heb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hec: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hf2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hf8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h116: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h11c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h122: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h128: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h12e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3a)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h134: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h135: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h138: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h139: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h13e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h13f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h144: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h145: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h14b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h151: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h157: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h15d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h163: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h169: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h16a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h16d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h16e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h173: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h174: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h179: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h17a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h180: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h186: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h18c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h192: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h198: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h19e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h19f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1a2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1a3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1a8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1a9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1ae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1af: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1b5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1bb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1c1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1c7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1cd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1d3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1d4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1d7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1d8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1dd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1de: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1e3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1e4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1ea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1f0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1f6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1fc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h202: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h20)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h4a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h50: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h56: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h62: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h68: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h6e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h74: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h7a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h7f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h85: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h8a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h8b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h91: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h97: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h9d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'haf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hba: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hbf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hcc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hde: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'he9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'heb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hec: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hfe: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h104: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h110: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h116: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h11c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h122: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h128: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h12e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h39)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3a)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h134: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h135: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h138: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h139: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h13e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h13f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h144: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h145: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h14b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h151: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h157: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h163: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h169: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h16a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h16d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h16e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h173: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h174: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h179: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h17a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h180: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h186: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h18c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h192: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h198: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h19e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h19f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1ae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1af: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1bb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1cd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1dd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1de: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1e3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ea: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1fc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h202: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						10'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						10'h207: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp22[14:0] );

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp255[14:0] );

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp470[14:0] );

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp685[14:0] );

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp900[14:0] );

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1115[14:0] );

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1330[14:0] );

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1545[14:0] );

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1760[14:0] );

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1978[14:0] );

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2193[14:0] );

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2408[14:0] );

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2623[14:0] );

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2838[14:0] );

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3053[14:0] );

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3268[14:0] );

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3483[14:0] );

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3701[14:0] );

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp3916[14:0] );

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4131[14:0] );

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4346[14:0] );

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4561[14:0] );

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4776[14:0] );

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp4991[14:0] );

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp5206[14:0] );

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp5424[14:0] );

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp5639[14:0] );

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp5854[14:0] );

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6069[14:0] );

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6284[14:0] );

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6499[14:0] );

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6714[14:0] );

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp6929[14:0] );

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11463[14:0] );

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11540[14:0] );

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11636[14:0] );

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11732[14:0] );

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11828[14:0] );

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11924[14:0] );

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12020[14:0] );

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12116[14:0] );

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12215[14:0] );

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12292[14:0] );

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12388[14:0] );

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12484[14:0] );

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12580[14:0] );

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12676[14:0] );

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12772[14:0] );

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12868[14:0] );

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12967[14:0] );

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13044[14:0] );

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13140[14:0] );

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13236[14:0] );

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13332[14:0] );

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13428[14:0] );

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13524[14:0] );

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13620[14:0] );

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13719[14:0] );

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13796[14:0] );

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13892[14:0] );

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13988[14:0] );

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp14084[14:0] );

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp14180[14:0] );

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp14276[14:0] );

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp14372[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11466;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11543;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11639;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11735;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11831;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp11927;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12023;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12119;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12218;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12295;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12391;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12487;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12583;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12679;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12775;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12871;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12970;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13047;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13143;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13239;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13335;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13431;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13527;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13623;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13722;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13799;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13895;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp13991;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp14087;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp14183;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp14279;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp14375;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h207: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp27[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h207: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp32[14:0] );

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp239[14:0] );

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp454[14:0] );

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp669[14:0] );

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp884[14:0] );

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1099[14:0] );

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1314[14:0] );

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1529[14:0] );

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1744[14:0] );

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1962[14:0] );

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2177[14:0] );

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2392[14:0] );

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2607[14:0] );

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2822[14:0] );

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3037[14:0] );

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3252[14:0] );

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3467[14:0] );

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3685[14:0] );

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3900[14:0] );

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4115[14:0] );

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4330[14:0] );

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4545[14:0] );

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4760[14:0] );

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4975[14:0] );

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5190[14:0] );

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5408[14:0] );

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5623[14:0] );

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5838[14:0] );

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6053[14:0] );

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6268[14:0] );

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6483[14:0] );

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6698[14:0] );

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6913[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp41[14:0] );

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp247[14:0] );

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp462[14:0] );

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp677[14:0] );

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp892[14:0] );

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1107[14:0] );

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1322[14:0] );

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1537[14:0] );

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1752[14:0] );

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1970[14:0] );

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2185[14:0] );

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2400[14:0] );

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2615[14:0] );

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2830[14:0] );

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3045[14:0] );

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3260[14:0] );

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3475[14:0] );

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3693[14:0] );

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3908[14:0] );

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4123[14:0] );

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4338[14:0] );

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4553[14:0] );

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4768[14:0] );

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4983[14:0] );

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5198[14:0] );

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5416[14:0] );

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5631[14:0] );

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5846[14:0] );

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6061[14:0] );

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6276[14:0] );

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6491[14:0] );

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6706[14:0] );

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6921[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_fld_V_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp14;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h11: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp229;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h46: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp1952;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h7b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp3675;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'hb0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp5398;

									end
								end

							endcase
						end

						10'heb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp7121;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_36 <= w_sys_tmp7204;

									end
								end

							endcase
						end

						10'hf1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp7205;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_36 <= w_sys_tmp7288;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp7289;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_36 <= w_sys_tmp7372;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp7373;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_36 <= w_sys_tmp7456;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp11452;

									end
								end

							endcase
						end

						10'h135: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp11456;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp12204;

									end
								end

							endcase
						end

						10'h16a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp12208;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp12956;

									end
								end

							endcase
						end

						10'h19f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp12960;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp13708;

									end
								end

							endcase
						end

						10'h1d4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_36 <= w_sys_tmp13712;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp48;

									end
								end

							endcase
						end

						10'h14: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp263;

									end
								end

							endcase
						end

						10'h1a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp444;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp478;

									end
								end

							endcase
						end

						10'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp659;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp693;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp874;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp908;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp1089;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp1123;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp1304;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp1338;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp1519;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp1553;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp1734;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp1768;

									end
								end

							endcase
						end

						10'h49: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp1986;

									end
								end

							endcase
						end

						10'h4f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp2167;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp2201;

									end
								end

							endcase
						end

						10'h55: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp2382;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp2416;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp2597;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp2631;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp2812;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp2846;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp3027;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp3061;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp3242;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp3276;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp3457;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp3491;

									end
								end

							endcase
						end

						10'h7e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp3709;

									end
								end

							endcase
						end

						10'h84: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp3890;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp3924;

									end
								end

							endcase
						end

						10'h8a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp4105;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp4139;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp4320;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp4354;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp4535;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp4569;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp4750;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp4784;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp4965;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp4999;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp5180;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp5214;

									end
								end

							endcase
						end

						10'hb3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp5432;

									end
								end

							endcase
						end

						10'hb9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp5613;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp5647;

									end
								end

							endcase
						end

						10'hbf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp5828;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp5862;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp6043;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp6077;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp6258;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp6292;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp6473;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp6507;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp6688;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp6722;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp6903;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp6937;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_37 <= w_sys_tmp7530;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp7957;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_37 <= w_sys_tmp8031;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp8458;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_37 <= w_sys_tmp8532;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp8959;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_37 <= w_sys_tmp9033;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp9460;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_37 <= w_sys_tmp9534;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp9961;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_37 <= w_sys_tmp10035;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp10462;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_37 <= w_sys_tmp10536;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp10963;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_37 <= w_sys_tmp11037;

									end
								end

							endcase
						end

						10'h138: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp11457;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp11471;

									end
								end

							endcase
						end

						10'h13e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp11532;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp11549;

									end
								end

							endcase
						end

						10'h144: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp11628;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp11645;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp11724;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp11741;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp11820;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp11837;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp11916;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp11933;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12012;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp12029;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12108;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp12125;

									end
								end

							endcase
						end

						10'h16d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12209;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp12223;

									end
								end

							endcase
						end

						10'h173: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12284;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp12301;

									end
								end

							endcase
						end

						10'h179: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12380;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp12397;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12476;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp12493;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12572;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp12589;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12668;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp12685;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12764;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp12781;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12860;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp12877;

									end
								end

							endcase
						end

						10'h1a2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp12961;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp12975;

									end
								end

							endcase
						end

						10'h1a8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13036;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp13053;

									end
								end

							endcase
						end

						10'h1ae: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13132;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp13149;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13228;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp13245;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13324;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp13341;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13420;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp13437;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13516;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp13533;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13612;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp13629;

									end
								end

							endcase
						end

						10'h1d7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13713;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_37 <= w_sys_tmp13727;

									end
								end

							endcase
						end

						10'h1dd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13788;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp13805;

									end
								end

							endcase
						end

						10'h1e3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13884;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp13901;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp13980;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp13997;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp14076;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp14093;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp14172;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp14189;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp14268;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp14285;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_37 <= w_sys_tmp14364;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_37 <= w_sys_tmp14381;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_38 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'he5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_38 <= w_sys_tmp7120;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_mx_39 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_my_40 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dt_41 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dx_42 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_dy_43 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r1_44 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r2_45 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r3_46 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_r4_47 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h10) || (r_sys_run_step==6'h11)) begin
										r_run_YY_48 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h14)) begin
										r_run_YY_48 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_kx_49 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_ky_50 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_nlast_51 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp11537;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp11633;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp11729;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp11825;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp11921;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp12017;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp12113;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp12289;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp12385;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp12481;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp12577;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp12673;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp12769;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp12865;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp13041;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp13137;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp13233;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp13329;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp13425;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp13521;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp13617;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp13793;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp13889;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp13985;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp14081;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp14177;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp14273;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_52 <= w_sys_tmp14369;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_53 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_53 <= w_sys_tmp45;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_54 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h18) || (r_sys_run_step==6'h1a) || (6'h1c<=r_sys_run_step && r_sys_run_step<=6'h20)) begin
										r_run_copy1_j_54 <= w_sys_tmp46;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_55 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_55 <= w_sys_tmp47;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_56 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_56 <= w_sys_tmp258;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_57 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_57 <= w_sys_tmp259;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_58 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_58 <= w_sys_tmp260;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_59 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_59 <= w_sys_tmp261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_60 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_60 <= w_sys_tmp262;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_61 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_61 <= w_sys_tmp473;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_62 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_62 <= w_sys_tmp474;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_63 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_63 <= w_sys_tmp475;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_64 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_64 <= w_sys_tmp476;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_65 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_65 <= w_sys_tmp477;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_66 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_66 <= w_sys_tmp688;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_67 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_67 <= w_sys_tmp689;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_68 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_68 <= w_sys_tmp690;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_69 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_69 <= w_sys_tmp691;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h20: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_70 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_70 <= w_sys_tmp692;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_71 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_71 <= w_sys_tmp903;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_72 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_72 <= w_sys_tmp904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_73 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_73 <= w_sys_tmp905;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_74 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_74 <= w_sys_tmp906;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_75 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_75 <= w_sys_tmp907;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_76 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_76 <= w_sys_tmp1118;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_77 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_77 <= w_sys_tmp1119;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_78 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_78 <= w_sys_tmp1120;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_79 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_79 <= w_sys_tmp1121;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_80 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_80 <= w_sys_tmp1122;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h32: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_81 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_81 <= w_sys_tmp1333;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h32: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_82 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_82 <= w_sys_tmp1334;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h32: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_83 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_83 <= w_sys_tmp1335;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h32: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_84 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_84 <= w_sys_tmp1336;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h32: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_85 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_85 <= w_sys_tmp1337;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h38: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_86 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_86 <= w_sys_tmp1548;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h38: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_87 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_87 <= w_sys_tmp1549;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h38: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_88 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_88 <= w_sys_tmp1550;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h38: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_89 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_89 <= w_sys_tmp1551;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h38: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_90 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_90 <= w_sys_tmp1552;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_91 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_91 <= w_sys_tmp1763;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_92 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_92 <= w_sys_tmp1764;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_93 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_93 <= w_sys_tmp1765;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_94 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_94 <= w_sys_tmp1766;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_95 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_95 <= w_sys_tmp1767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h49: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_96 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_96 <= w_sys_tmp1981;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h49: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_97 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_97 <= w_sys_tmp1982;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h49: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_98 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_98 <= w_sys_tmp1983;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h49: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_99 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_99 <= w_sys_tmp1984;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h49: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_100 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_100 <= w_sys_tmp1985;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_101 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_101 <= w_sys_tmp2196;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_102 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_102 <= w_sys_tmp2197;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_103 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_103 <= w_sys_tmp2198;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_104 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_104 <= w_sys_tmp2199;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_105 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_105 <= w_sys_tmp2200;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h55: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_106 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_106 <= w_sys_tmp2411;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h55: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_107 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_107 <= w_sys_tmp2412;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h55: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_108 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_108 <= w_sys_tmp2413;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h55: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_109 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_109 <= w_sys_tmp2414;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h55: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_110 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_110 <= w_sys_tmp2415;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_111 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_111 <= w_sys_tmp2626;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_112 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_112 <= w_sys_tmp2627;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_113 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_113 <= w_sys_tmp2628;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_114 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_114 <= w_sys_tmp2629;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_115 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_115 <= w_sys_tmp2630;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h61: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_116 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_116 <= w_sys_tmp2841;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h61: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_117 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_117 <= w_sys_tmp2842;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h61: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_118 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_118 <= w_sys_tmp2843;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h61: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_119 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_119 <= w_sys_tmp2844;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h61: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_120 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_120 <= w_sys_tmp2845;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h67: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_121 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_121 <= w_sys_tmp3056;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h67: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_122 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_122 <= w_sys_tmp3057;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h67: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_123 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_123 <= w_sys_tmp3058;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h67: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_124 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_124 <= w_sys_tmp3059;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h67: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_125 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_125 <= w_sys_tmp3060;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_126 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_126 <= w_sys_tmp3271;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_127 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_127 <= w_sys_tmp3272;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_128 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_128 <= w_sys_tmp3273;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_129 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_129 <= w_sys_tmp3274;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_130 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_130 <= w_sys_tmp3275;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h73: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_131 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_131 <= w_sys_tmp3486;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h73: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_132 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_132 <= w_sys_tmp3487;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h73: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_133 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_133 <= w_sys_tmp3488;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h73: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_134 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_134 <= w_sys_tmp3489;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h73: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_135 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_135 <= w_sys_tmp3490;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_136 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_136 <= w_sys_tmp3704;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_137 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_137 <= w_sys_tmp3705;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_138 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_138 <= w_sys_tmp3706;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_139 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_139 <= w_sys_tmp3707;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_140 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_140 <= w_sys_tmp3708;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h84: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_141 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_141 <= w_sys_tmp3919;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h84: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_142 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_142 <= w_sys_tmp3920;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h84: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_143 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_143 <= w_sys_tmp3921;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h84: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_144 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_144 <= w_sys_tmp3922;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h84: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_145 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_145 <= w_sys_tmp3923;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_146 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_146 <= w_sys_tmp4134;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_147 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_147 <= w_sys_tmp4135;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_148 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_148 <= w_sys_tmp4136;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_149 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_149 <= w_sys_tmp4137;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_150 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_150 <= w_sys_tmp4138;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h90: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_151 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_151 <= w_sys_tmp4349;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h90: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_152 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_152 <= w_sys_tmp4350;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h90: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_153 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_153 <= w_sys_tmp4351;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h90: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_154 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_154 <= w_sys_tmp4352;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h90: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_155 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_155 <= w_sys_tmp4353;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h96: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_156 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_156 <= w_sys_tmp4564;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h96: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_157 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_157 <= w_sys_tmp4565;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h96: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_158 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_158 <= w_sys_tmp4566;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h96: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_159 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_159 <= w_sys_tmp4567;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h96: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_160 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_160 <= w_sys_tmp4568;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_161 <= r_run_j_37;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_161 <= w_sys_tmp4779;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_162 <= r_run_j_37;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_162 <= w_sys_tmp4780;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_163 <= r_run_j_37;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_163 <= w_sys_tmp4781;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_164 <= r_run_j_37;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_164 <= w_sys_tmp4782;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_165 <= r_run_j_37;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_165 <= w_sys_tmp4783;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_166 <= r_run_j_37;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_166 <= w_sys_tmp4994;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_167 <= r_run_j_37;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_167 <= w_sys_tmp4995;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_168 <= r_run_j_37;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_168 <= w_sys_tmp4996;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_169 <= r_run_j_37;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_169 <= w_sys_tmp4997;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_170 <= r_run_j_37;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_170 <= w_sys_tmp4998;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_171 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_171 <= w_sys_tmp5209;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_172 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_172 <= w_sys_tmp5210;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_173 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_173 <= w_sys_tmp5211;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_174 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_174 <= w_sys_tmp5212;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_175 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_175 <= w_sys_tmp5213;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_176 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_176 <= w_sys_tmp5427;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_177 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_177 <= w_sys_tmp5428;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_178 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_178 <= w_sys_tmp5429;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_179 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_179 <= w_sys_tmp5430;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_180 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_180 <= w_sys_tmp5431;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_181 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_181 <= w_sys_tmp5642;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_182 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_182 <= w_sys_tmp5643;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_183 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_183 <= w_sys_tmp5644;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_184 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_184 <= w_sys_tmp5645;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_185 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_185 <= w_sys_tmp5646;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_186 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_186 <= w_sys_tmp5857;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_187 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_187 <= w_sys_tmp5858;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_188 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_188 <= w_sys_tmp5859;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_189 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_189 <= w_sys_tmp5860;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbf: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_190 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_190 <= w_sys_tmp5861;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_191 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_191 <= w_sys_tmp6072;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_192 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_192 <= w_sys_tmp6073;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_193 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_193 <= w_sys_tmp6074;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_194 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_194 <= w_sys_tmp6075;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_195 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_195 <= w_sys_tmp6076;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcb: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_196 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_196 <= w_sys_tmp6287;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcb: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_197 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_197 <= w_sys_tmp6288;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcb: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_198 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_198 <= w_sys_tmp6289;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcb: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_199 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_199 <= w_sys_tmp6290;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcb: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_200 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_200 <= w_sys_tmp6291;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd1: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_201 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_201 <= w_sys_tmp6502;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd1: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_202 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_202 <= w_sys_tmp6503;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd1: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_203 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_203 <= w_sys_tmp6504;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd1: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_204 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_204 <= w_sys_tmp6505;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd1: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_205 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_205 <= w_sys_tmp6506;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd7: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_206 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_206 <= w_sys_tmp6717;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd7: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_207 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_207 <= w_sys_tmp6718;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd7: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_208 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_208 <= w_sys_tmp6719;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd7: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_209 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_209 <= w_sys_tmp6720;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd7: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_210 <= r_run_j_37;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_210 <= w_sys_tmp6721;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_211 <= r_run_j_37;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_211 <= w_sys_tmp6932;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_212 <= r_run_j_37;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_212 <= w_sys_tmp6933;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_213 <= r_run_j_37;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy2_j_213 <= w_sys_tmp6934;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_214 <= r_run_j_37;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy3_j_214 <= w_sys_tmp6935;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_215 <= r_run_j_37;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy4_j_215 <= w_sys_tmp6936;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_216 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_216 <= w_sys_tmp7519;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_217 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_217 <= w_sys_tmp7520;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_218 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_218 <= w_sys_tmp7521;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_219 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_219 <= w_sys_tmp7522;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_220 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_220 <= w_sys_tmp7523;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_221 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_221 <= w_sys_tmp7524;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_222 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_222 <= w_sys_tmp7525;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_223 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_223 <= w_sys_tmp7526;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_224 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_224 <= w_sys_tmp7527;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_225 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_225 <= w_sys_tmp7528;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_226 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_226 <= w_sys_tmp7529;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_227 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_227 <= w_sys_tmp8020;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_228 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_228 <= w_sys_tmp8021;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_229 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_229 <= w_sys_tmp8022;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_230 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_230 <= w_sys_tmp8023;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_231 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_231 <= w_sys_tmp8024;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_232 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_232 <= w_sys_tmp8025;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_233 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_233 <= w_sys_tmp8026;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_234 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_234 <= w_sys_tmp8027;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_235 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_235 <= w_sys_tmp8028;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_236 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_236 <= w_sys_tmp8029;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_237 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_237 <= w_sys_tmp8030;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_238 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_238 <= w_sys_tmp8521;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_239 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_239 <= w_sys_tmp8522;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_240 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_240 <= w_sys_tmp8523;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_241 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_241 <= w_sys_tmp8524;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_242 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_242 <= w_sys_tmp8525;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_243 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_243 <= w_sys_tmp8526;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_244 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_244 <= w_sys_tmp8527;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_245 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_245 <= w_sys_tmp8528;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_246 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_246 <= w_sys_tmp8529;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_247 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_247 <= w_sys_tmp8530;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_248 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_248 <= w_sys_tmp8531;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_249 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_249 <= w_sys_tmp9022;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_250 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_250 <= w_sys_tmp9023;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_251 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_251 <= w_sys_tmp9024;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_252 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_252 <= w_sys_tmp9025;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_253 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_253 <= w_sys_tmp9026;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_254 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_254 <= w_sys_tmp9027;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_255 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_255 <= w_sys_tmp9028;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_256 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_256 <= w_sys_tmp9029;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_257 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_257 <= w_sys_tmp9030;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_258 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_258 <= w_sys_tmp9031;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_259 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_259 <= w_sys_tmp9032;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_260 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_260 <= w_sys_tmp9523;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_261 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_261 <= w_sys_tmp9524;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_262 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_262 <= w_sys_tmp9525;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_263 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_263 <= w_sys_tmp9526;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_264 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_264 <= w_sys_tmp9527;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_265 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_265 <= w_sys_tmp9528;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_266 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_266 <= w_sys_tmp9529;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_267 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_267 <= w_sys_tmp9530;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_268 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_268 <= w_sys_tmp9531;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_269 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_269 <= w_sys_tmp9532;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_270 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_270 <= w_sys_tmp9533;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_271 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_271 <= w_sys_tmp10024;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_272 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_272 <= w_sys_tmp10025;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_273 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_273 <= w_sys_tmp10026;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_274 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_274 <= w_sys_tmp10027;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_275 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_275 <= w_sys_tmp10028;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_276 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_276 <= w_sys_tmp10029;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_277 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_277 <= w_sys_tmp10030;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_278 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_278 <= w_sys_tmp10031;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_279 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_279 <= w_sys_tmp10032;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_280 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_280 <= w_sys_tmp10033;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_281 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_281 <= w_sys_tmp10034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_282 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_282 <= w_sys_tmp10525;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_283 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_283 <= w_sys_tmp10526;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_284 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_284 <= w_sys_tmp10527;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_285 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_285 <= w_sys_tmp10528;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_286 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_286 <= w_sys_tmp10529;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_287 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_287 <= w_sys_tmp10530;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_288 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_288 <= w_sys_tmp10531;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_289 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_289 <= w_sys_tmp10532;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_290 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_290 <= w_sys_tmp10533;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_291 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_291 <= w_sys_tmp10534;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_292 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_292 <= w_sys_tmp10535;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_293 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_293 <= w_sys_tmp11026;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_294 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'he)) begin
										r_run_copy1_j_294 <= w_sys_tmp11027;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_295 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_run_copy2_j_295 <= w_sys_tmp11028;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_296 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_296 <= w_sys_tmp11029;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_297 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_297 <= w_sys_tmp11030;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_298 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_298 <= w_sys_tmp11031;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_299 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy6_j_299 <= w_sys_tmp11032;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_300 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_300 <= w_sys_tmp11033;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_301 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_301 <= w_sys_tmp11034;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_302 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_302 <= w_sys_tmp11035;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_303 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_303 <= w_sys_tmp11036;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h138: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_304 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_304 <= w_sys_tmp11470;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_305 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_305 <= w_sys_tmp11547;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13e: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_306 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_306 <= w_sys_tmp11548;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h144: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_307 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_307 <= w_sys_tmp11643;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h144: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_308 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_308 <= w_sys_tmp11644;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_309 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_309 <= w_sys_tmp11739;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14a: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_310 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_310 <= w_sys_tmp11740;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h150: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_311 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_311 <= w_sys_tmp11835;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h150: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_312 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_312 <= w_sys_tmp11836;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h156: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_313 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_313 <= w_sys_tmp11931;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h156: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_314 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_314 <= w_sys_tmp11932;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h15c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_315 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_315 <= w_sys_tmp12027;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h15c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_316 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_316 <= w_sys_tmp12028;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h162: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_317 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_317 <= w_sys_tmp12123;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h162: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_318 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_318 <= w_sys_tmp12124;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h16d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_319 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_319 <= w_sys_tmp12222;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h173: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_320 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_320 <= w_sys_tmp12299;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h173: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_321 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_321 <= w_sys_tmp12300;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h179: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_322 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_322 <= w_sys_tmp12395;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h179: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_323 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_323 <= w_sys_tmp12396;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h17f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_324 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_324 <= w_sys_tmp12491;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h17f: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_325 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_325 <= w_sys_tmp12492;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h185: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_326 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_326 <= w_sys_tmp12587;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h185: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_327 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_327 <= w_sys_tmp12588;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_328 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_328 <= w_sys_tmp12683;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18b: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_329 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_329 <= w_sys_tmp12684;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h191: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_330 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_330 <= w_sys_tmp12779;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h191: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_331 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_331 <= w_sys_tmp12780;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h197: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_332 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_332 <= w_sys_tmp12875;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h197: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_333 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_333 <= w_sys_tmp12876;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a2: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_334 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_334 <= w_sys_tmp12974;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_335 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_335 <= w_sys_tmp13051;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a8: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_336 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_336 <= w_sys_tmp13052;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ae: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_337 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_337 <= w_sys_tmp13147;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ae: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_338 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_338 <= w_sys_tmp13148;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1b4: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_339 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_339 <= w_sys_tmp13243;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1b4: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_340 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_340 <= w_sys_tmp13244;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ba: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_341 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_341 <= w_sys_tmp13339;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ba: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_342 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_342 <= w_sys_tmp13340;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_343 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_343 <= w_sys_tmp13435;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c0: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_344 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_344 <= w_sys_tmp13436;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_345 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_345 <= w_sys_tmp13531;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c6: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_346 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_346 <= w_sys_tmp13532;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1cc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_347 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_347 <= w_sys_tmp13627;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1cc: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_348 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_348 <= w_sys_tmp13628;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1d7: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_349 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_349 <= w_sys_tmp13726;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1dd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_350 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_350 <= w_sys_tmp13803;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1dd: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_351 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_351 <= w_sys_tmp13804;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_352 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_352 <= w_sys_tmp13899;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e3: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_353 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_353 <= w_sys_tmp13900;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_354 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_354 <= w_sys_tmp13995;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_355 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_355 <= w_sys_tmp13996;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_356 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_356 <= w_sys_tmp14091;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ef: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_357 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_357 <= w_sys_tmp14092;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1f5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_358 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_358 <= w_sys_tmp14187;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1f5: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_359 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_359 <= w_sys_tmp14188;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1fb: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_360 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_360 <= w_sys_tmp14283;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1fb: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_361 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_361 <= w_sys_tmp14284;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h201: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_362 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_362 <= w_sys_tmp14379;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h201: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_363 <= r_run_j_37;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_363 <= w_sys_tmp14380;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp4342[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_T_datain <= w_sys_tmp4345;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub19_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp4334[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_V_datain <= w_sys_tmp4337;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub19_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp4326[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_U_datain <= w_sys_tmp4329;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub19_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hf)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp7295[14:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp7307[14:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp7301[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp7298[14:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp9018[14:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp9004[14:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp8994[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp8989[14:0] );

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp13240[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub19_result_datain <= w_sys_tmp7325;

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub19_result_datain <= r_sys_tmp4_float;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub19_result_datain <= w_sys_tmp8969;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub19_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'hf)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub19_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub19_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub19_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp2834[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_T_datain <= w_sys_tmp2837;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub12_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp2826[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_V_datain <= w_sys_tmp2829;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub12_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp2818[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_U_datain <= w_sys_tmp2821;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub12_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp7223[14:0] );

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp7217[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp7214[14:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp7211[14:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp9476[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp9471[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp9486[14:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp9500[14:0] );

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12584[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub12_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub12_result_datain <= w_sys_tmp7252;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub12_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub12_result_datain <= w_sys_tmp9518;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub12_result_datain <= w_sys_tmp9480;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp2619[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_T_datain <= w_sys_tmp2622;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub11_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp2611[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_V_datain <= w_sys_tmp2614;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub11_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp2603[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_U_datain <= w_sys_tmp2606;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub11_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp7223[14:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp7217[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp7214[14:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp7211[14:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp8970[14:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp8975[14:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp8999[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp8985[14:0] );

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12488[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub11_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub11_result_datain <= w_sys_tmp7241;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub11_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub11_result_datain <= w_sys_tmp8979;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_datain <= w_sys_tmp9017;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hf)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp3264[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_T_datain <= w_sys_tmp3267;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub14_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp3256[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_V_datain <= w_sys_tmp3259;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub14_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp3248[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_U_datain <= w_sys_tmp3251;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub14_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp7223[14:0] );

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp7217[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp7214[14:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp7211[14:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp10502[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp10473[14:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp10478[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp10488[14:0] );

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12776[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub14_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub14_result_datain <= w_sys_tmp7274;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub14_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub14_result_datain <= w_sys_tmp10482;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub14_result_datain <= w_sys_tmp10520;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp3049[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_T_datain <= w_sys_tmp3052;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub13_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp3041[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_V_datain <= w_sys_tmp3044;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub13_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp3033[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_U_datain <= w_sys_tmp3036;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub13_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp7223[14:0] );

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp7217[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp7214[14:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp7211[14:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp10001[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp9972[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp9987[14:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp9977[14:0] );

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12680[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h15)) begin
										r_sub13_result_datain <= w_sys_tmp7263;

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub13_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub13_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub13_result_datain <= w_sys_tmp9981;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_datain <= w_sys_tmp10019;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp3697[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_T_datain <= w_sys_tmp3700;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub16_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp3689[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_V_datain <= w_sys_tmp3692;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub16_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp3681[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_U_datain <= w_sys_tmp3684;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub16_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp7295[14:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp7304[14:0] );

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp7501[14:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp7515[14:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp7491[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp7486[14:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp11022[14:0] );

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12971[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub16_result_datain <= w_sys_tmp7297;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub16_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub16_result_datain <= w_sys_tmp7466;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub16_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub16_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub16_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp3479[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_T_datain <= w_sys_tmp3482;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub15_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp3471[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_V_datain <= w_sys_tmp3474;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub15_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp3463[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_U_datain <= w_sys_tmp3466;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub15_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp7217[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp7214[14:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp10974[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp10989[14:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp11003[14:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp10979[14:0] );

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12872[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub15_result_datain <= w_sys_tmp7285;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_datain <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub15_result_datain <= w_sys_tmp10983;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp4127[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_T_datain <= w_sys_tmp4130;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub18_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp4119[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_V_datain <= w_sys_tmp4122;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub18_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp4111[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_U_datain <= w_sys_tmp4114;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub18_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp7295[14:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp7307[14:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp7301[14:0] );

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp8503[14:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp8517[14:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp8493[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp8488[14:0] );

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp13144[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub18_result_datain <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub18_result_datain <= w_sys_tmp7297;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub18_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub18_result_datain <= w_sys_tmp8468;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub18_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub18_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub18_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp3912[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_T_datain <= w_sys_tmp3915;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub17_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp3904[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_V_datain <= w_sys_tmp3907;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub17_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp3896[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_U_datain <= w_sys_tmp3899;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub17_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp7295[14:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp7307[14:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp7301[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp7298[14:0] );

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp7992[14:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp8016[14:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp8002[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp7987[14:0] );

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp13048[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub17_result_datain <= w_sys_tmp7303;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub17_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub17_result_datain <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub17_result_datain <= w_sys_tmp7967;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub17_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub17_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub17_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp4557[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_T_datain <= w_sys_tmp4560;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub20_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp4549[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_V_datain <= w_sys_tmp4552;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub20_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp4541[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_U_datain <= w_sys_tmp4544;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub20_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h13)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp7295[14:0] );

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp7307[14:0] );

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp7301[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp7298[14:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp9519[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp9490[14:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp9495[14:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp9505[14:0] );

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13336[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub20_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub20_result_datain <= w_sys_tmp7336;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub20_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub20_result_datain <= w_sys_tmp9470;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub20_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub20_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub20_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp4772[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_T_datain <= w_sys_tmp4775;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub21_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp4764[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_V_datain <= w_sys_tmp4767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub21_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp4756[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_U_datain <= w_sys_tmp4759;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub21_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h17)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp7295[14:0] );

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp7307[14:0] );

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp7301[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp7298[14:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp9996[14:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp10006[14:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp10020[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp9991[14:0] );

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13432[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub21_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub21_result_datain <= w_sys_tmp7347;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub21_result_datain <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub21_result_datain <= w_sys_tmp9971;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub21_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub21_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub21_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_T_addr <= $signed( w_sys_tmp6280[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_T_datain <= w_sys_tmp6283;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub28_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_V_addr <= $signed( w_sys_tmp6272[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_V_datain <= w_sys_tmp6275;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub28_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_U_addr <= $signed( w_sys_tmp6264[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_U_datain <= w_sys_tmp6267;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub28_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp7385[14:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp7379[14:0] );

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp7391[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp7382[14:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp9509[14:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp9514[14:0] );

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp14088[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub28_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub28_result_datain <= w_sys_tmp7420;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub28_result_datain <= w_sys_tmp9518;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub28_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub28_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub28_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_T_addr <= $signed( w_sys_tmp6495[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_T_datain <= w_sys_tmp6498;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub29_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_V_addr <= $signed( w_sys_tmp6487[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_V_datain <= w_sys_tmp6490;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub29_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_U_addr <= $signed( w_sys_tmp6479[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_U_datain <= w_sys_tmp6482;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub29_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h15)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp7385[14:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp7379[14:0] );

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp7391[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp7382[14:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp10015[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp10010[14:0] );

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp14184[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h15)) begin
										r_sub29_result_datain <= w_sys_tmp7431;

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub29_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub29_result_datain <= w_sys_tmp10019;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub29_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub29_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub29_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_T_addr <= $signed( w_sys_tmp5850[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_T_datain <= w_sys_tmp5853;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub26_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_V_addr <= $signed( w_sys_tmp5842[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_V_datain <= w_sys_tmp5845;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub26_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_U_addr <= $signed( w_sys_tmp5834[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_U_datain <= w_sys_tmp5837;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub26_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp7385[14:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp7379[14:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp7391[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp7382[14:0] );

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp8507[14:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp8512[14:0] );

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp13896[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub26_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub26_result_datain <= w_sys_tmp7381;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub26_result_datain <= w_sys_tmp8516;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub26_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub26_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub26_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp2189[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_T_datain <= w_sys_tmp2192;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub09_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp2181[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_V_datain <= w_sys_tmp2184;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub09_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp2173[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_U_datain <= w_sys_tmp2176;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub09_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp7223[14:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp7217[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp7214[14:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp7211[14:0] );

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp7973[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp7968[14:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp7997[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp7983[14:0] );

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp12296[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub09_result_datain <= w_sys_tmp7219;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub09_result_datain <= w_sys_tmp7977;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_datain <= w_sys_tmp8015;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_T_addr <= $signed( w_sys_tmp6065[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_T_datain <= w_sys_tmp6068;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub27_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_V_addr <= $signed( w_sys_tmp6057[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_V_datain <= w_sys_tmp6060;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub27_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_U_addr <= $signed( w_sys_tmp6049[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_U_datain <= w_sys_tmp6052;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub27_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp7385[14:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp7379[14:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp7391[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp7382[14:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp9008[14:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp9013[14:0] );

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp13992[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub27_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub27_result_datain <= w_sys_tmp7409;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub27_result_datain <= w_sys_tmp9017;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hf)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub27_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub27_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub27_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp1974[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_T_datain <= w_sys_tmp1977;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub08_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1966[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_V_datain <= w_sys_tmp1969;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub08_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1958[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_U_datain <= w_sys_tmp1961;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub08_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp7220[14:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp7211[14:0] );

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp7482[14:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp7472[14:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp7496[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp7467[14:0] );

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp12219[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub08_result_datain <= w_sys_tmp7213;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub08_result_datain <= w_sys_tmp7476;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub08_result_datain <= w_sys_tmp7514;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub08_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp5420[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_T_datain <= w_sys_tmp5423;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub24_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp5412[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_V_datain <= w_sys_tmp5415;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub24_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp5404[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_U_datain <= w_sys_tmp5407;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub24_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp7379[14:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp7388[14:0] );

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp7510[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp7505[14:0] );

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13723[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub24_result_datain <= w_sys_tmp7381;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub24_result_datain <= w_sys_tmp7514;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub24_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub24_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub24_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_T_addr <= $signed( w_sys_tmp5635[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_T_datain <= w_sys_tmp5638;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub25_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_V_addr <= $signed( w_sys_tmp5627[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_V_datain <= w_sys_tmp5630;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub25_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_U_addr <= $signed( w_sys_tmp5619[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_U_datain <= w_sys_tmp5622;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub25_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp7385[14:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp7379[14:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp7391[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp7382[14:0] );

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp8006[14:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp8011[14:0] );

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp13800[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub25_result_datain <= w_sys_tmp7387;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub25_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub25_result_datain <= w_sys_tmp8015;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub25_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub25_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub25_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp4987[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_T_datain <= w_sys_tmp4990;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub22_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp4979[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_V_datain <= w_sys_tmp4982;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub22_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp4971[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_U_datain <= w_sys_tmp4974;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub22_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1b)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp7295[14:0] );

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp7307[14:0] );

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp7301[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp7298[14:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp10492[14:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp10507[14:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp10521[14:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp10497[14:0] );

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13528[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub22_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub22_result_datain <= w_sys_tmp7358;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub22_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub22_result_datain <= w_sys_tmp10472;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub22_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub22_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub22_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp5202[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_T_datain <= w_sys_tmp5205;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub23_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp5194[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_V_datain <= w_sys_tmp5197;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub23_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp5186[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_U_datain <= w_sys_tmp5189;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub23_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp7301[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp7298[14:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp11008[14:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp10998[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp10993[14:0] );

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13624[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub23_result_datain <= w_sys_tmp7369;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h32)) begin
										r_sub23_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h22)) begin
										r_sub23_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h2a)) begin
										r_sub23_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub23_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub23_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub23_result_datain <= w_sys_tmp10973;

									end
									else
									if((r_sys_run_step==6'h3a)) begin
										r_sub23_result_datain <= r_sys_tmp6_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub23_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub23_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub23_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp896[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_datain <= w_sys_tmp899;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub03_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp888[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_V_datain <= w_sys_tmp891;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub03_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp880[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_datain <= w_sys_tmp883;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub03_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp7133[14:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp7127[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp7130[14:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp7139[14:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp8980[14:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp8965[14:0] );

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11736[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub03_result_datain <= w_sys_tmp7157;

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub03_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub03_result_datain <= w_sys_tmp8969;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hf)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp681[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_datain <= w_sys_tmp684;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub02_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp673[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_V_datain <= w_sys_tmp676;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub02_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp665[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_datain <= w_sys_tmp668;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub02_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp7133[14:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp7127[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp7130[14:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp7139[14:0] );

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp8464[14:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp8479[14:0] );

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11640[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub02_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub02_result_datain <= w_sys_tmp7129;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub02_result_datain <= w_sys_tmp8468;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp466[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_datain <= w_sys_tmp469;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub01_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp458[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_V_datain <= w_sys_tmp461;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub01_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp450[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_datain <= w_sys_tmp453;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub01_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp7133[14:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp7127[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp7130[14:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp7139[14:0] );

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp7978[14:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp7963[14:0] );

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp11544[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub01_result_datain <= w_sys_tmp7135;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub01_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub01_result_datain <= w_sys_tmp7967;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp251[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_datain <= w_sys_tmp254;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub00_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp243[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_V_datain <= w_sys_tmp246;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub00_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp235[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_datain <= w_sys_tmp238;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub00_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp7127[14:0] );

									end
									else
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp7136[14:0] );

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp7477[14:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp7462[14:0] );

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp11467[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_datain <= w_sys_tmp7129;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_datain <= w_sys_tmp7466;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp1756[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_datain <= w_sys_tmp1759;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub07_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1748[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_V_datain <= w_sys_tmp1751;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub07_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1740[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_datain <= w_sys_tmp1743;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub07_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp7133[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp7130[14:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp10984[14:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp10969[14:0] );

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp12120[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub07_result_datain <= w_sys_tmp7201;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub07_result_datain <= w_sys_tmp10973;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp1541[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_datain <= w_sys_tmp1544;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub06_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1533[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_V_datain <= w_sys_tmp1536;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub06_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1525[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_datain <= w_sys_tmp1528;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub06_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h19)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp7133[14:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp7127[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp7130[14:0] );

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp7139[14:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp10483[14:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp10468[14:0] );

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp12024[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub06_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub06_result_datain <= w_sys_tmp7190;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub06_result_datain <= w_sys_tmp10472;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp1326[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_datain <= w_sys_tmp1329;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub05_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1318[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_V_datain <= w_sys_tmp1321;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub05_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1310[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_datain <= w_sys_tmp1313;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub05_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h15)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp7133[14:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp7127[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp7130[14:0] );

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp7139[14:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp9982[14:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp9967[14:0] );

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11928[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub05_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub05_result_datain <= w_sys_tmp7179;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub05_result_datain <= w_sys_tmp9971;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1111[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_datain <= w_sys_tmp1114;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub04_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1103[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_V_datain <= w_sys_tmp1106;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub04_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1095[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_datain <= w_sys_tmp1098;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub04_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp7133[14:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp7127[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp7130[14:0] );

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp7139[14:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp9466[14:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp9481[14:0] );

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11832[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub04_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub04_result_datain <= w_sys_tmp7168;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_datain <= w_sys_tmp9470;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp2404[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_T_datain <= w_sys_tmp2407;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub10_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp2396[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_V_datain <= w_sys_tmp2399;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub10_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp2388[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_U_datain <= w_sys_tmp2391;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub10_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp7223[14:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp7217[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp7214[14:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp7211[14:0] );

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp8474[14:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp8484[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp8469[14:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp8498[14:0] );

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12392[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub10_result_datain <= w_sys_tmp7213;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub10_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub10_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub10_result_datain <= w_sys_tmp8516;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub10_result_datain <= w_sys_tmp8478;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_T_addr <= $signed( w_sys_tmp6925[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_T_datain <= w_sys_tmp6928;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub31_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_V_addr <= $signed( w_sys_tmp6917[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_V_datain <= w_sys_tmp6920;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub31_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_U_addr <= $signed( w_sys_tmp6909[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_U_datain <= w_sys_tmp6912;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub31_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp7385[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp7382[14:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp11012[14:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'he)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp11017[14:0] );

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp14376[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub31_result_datain <= w_sys_tmp7453;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub31_result_datain <= w_sys_tmp11021;

									end
									else
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'he)) begin
										r_sub31_result_datain <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'hc)) begin
										r_sub31_result_datain <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'ha)) begin
										r_sub31_result_datain <= r_sys_tmp6_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub31_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'he)) begin
										r_sub31_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub31_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_T_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_T_addr <= $signed( w_sys_tmp6710[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_T_datain <= w_sys_tmp6713;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub30_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_V_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_V_addr <= $signed( w_sys_tmp6702[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_V_datain <= w_sys_tmp6705;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub30_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_U_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_U_addr <= $signed( w_sys_tmp6694[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_U_datain <= w_sys_tmp6697;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub30_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_result_addr <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h19)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp7385[14:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp7379[14:0] );

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp7391[14:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp7382[14:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp10516[14:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp10511[14:0] );

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp14280[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub30_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub30_result_datain <= w_sys_tmp7442;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub30_result_datain <= w_sys_tmp10520;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub30_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub30_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub30_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub27_result_dataout;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp0_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp0_float <= w_sub28_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sys_tmp0_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub29_result_dataout;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub20_result_dataout;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_tmp1_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h12) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h19)) begin
										r_sys_tmp2_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp2_float <= w_sub26_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sys_tmp2_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h17)) begin
										r_sys_tmp3_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub30_result_dataout;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp3_float <= w_sub27_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sys_tmp3_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h19)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==6'hc) || (r_sys_run_step==6'hd)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub20_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub28_result_dataout;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp4_float <= w_sub30_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'hb)) begin
										r_sys_tmp4_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp5_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub26_result_dataout;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp5_float <= w_sub25_result_dataout;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp5_float <= w_sub29_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h8)) begin
										r_sys_tmp5_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'hf)) begin
										r_sys_tmp6_float <= w_sub31_result_dataout;

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6)) begin
										r_sys_tmp6_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h131: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sys_tmp7_float <= w_sub16_result_dataout;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sys_tmp7_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
