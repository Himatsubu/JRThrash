/*
TimeStamp:	2016/12/23		13:32
*/


module NeuralNetJRT(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_threadTop_req,	
	output                o_threadTop_busy	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg         [31:0] r_ip_DivFloat_dividend_0;
	reg         [31:0] r_ip_DivFloat_divisor_0;
	wire        [31:0] w_ip_DivFloat_quotient_0;
	reg         [31:0] r_ip_CompareFloatLT_portA_0;
	reg         [31:0] r_ip_CompareFloatLT_portB_0;
	wire               w_ip_CompareFloatLT_result_0;
	reg         [31:0] r_ip_exp_i_0;
	wire        [31:0] w_ip_exp_result_0;
	reg                r_ip_exp_newData_0;
	reg         [31:0] r_ip_exp_i_1;
	wire        [31:0] w_ip_exp_result_1;
	reg                r_ip_exp_newData_1;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_threadTop_caller;
	reg                r_sys_threadTop_req;
	reg         [ 6:0] r_sys_threadTop_phase;
	reg         [ 1:0] r_sys_threadTop_stage;
	reg         [ 6:0] r_sys_threadTop_step;
	reg                r_sys_threadTop_busy;
	wire        [ 1:0] w_sys_threadTop_stage_p1;
	wire        [ 6:0] w_sys_threadTop_step_p1;
	reg  signed [31:0] r_fld_N_INPUT_0;
	reg  signed [31:0] r_fld_N_HIDDEN_1;
	reg  signed [31:0] r_fld_N_OUTPUT_2;
	wire signed [ 3:0] w_fld_w1_3_addr_0;
	wire        [31:0] w_fld_w1_3_datain_0;
	wire        [31:0] w_fld_w1_3_dataout_0;
	wire               w_fld_w1_3_r_w_0;
	wire               w_fld_w1_3_ce_0;
	reg  signed [ 3:0] r_fld_w1_3_addr_1;
	reg         [31:0] r_fld_w1_3_datain_1;
	wire        [31:0] w_fld_w1_3_dataout_1;
	reg                r_fld_w1_3_r_w_1;
	wire               w_fld_w1_3_ce_1;
	wire signed [ 2:0] w_fld_w2_4_addr_0;
	wire        [31:0] w_fld_w2_4_datain_0;
	wire        [31:0] w_fld_w2_4_dataout_0;
	wire               w_fld_w2_4_r_w_0;
	wire               w_fld_w2_4_ce_0;
	reg  signed [ 2:0] r_fld_w2_4_addr_1;
	reg         [31:0] r_fld_w2_4_datain_1;
	wire        [31:0] w_fld_w2_4_dataout_1;
	reg                r_fld_w2_4_r_w_1;
	wire               w_fld_w2_4_ce_1;
	wire signed        w_fld_input_5_addr_0;
	wire        [31:0] w_fld_input_5_datain_0;
	wire        [31:0] w_fld_input_5_dataout_0;
	wire               w_fld_input_5_r_w_0;
	wire               w_fld_input_5_ce_0;
	reg  signed        r_fld_input_5_addr_1;
	reg         [31:0] r_fld_input_5_datain_1;
	wire        [31:0] w_fld_input_5_dataout_1;
	reg                r_fld_input_5_r_w_1;
	wire               w_fld_input_5_ce_1;
	wire signed [ 2:0] w_fld_hidden_6_addr_0;
	wire        [31:0] w_fld_hidden_6_datain_0;
	wire        [31:0] w_fld_hidden_6_dataout_0;
	wire               w_fld_hidden_6_r_w_0;
	wire               w_fld_hidden_6_ce_0;
	reg  signed [ 2:0] r_fld_hidden_6_addr_1;
	reg         [31:0] r_fld_hidden_6_datain_1;
	wire        [31:0] w_fld_hidden_6_dataout_1;
	reg                r_fld_hidden_6_r_w_1;
	wire               w_fld_hidden_6_ce_1;
	wire signed        w_fld_output_7_addr_0;
	wire        [31:0] w_fld_output_7_datain_0;
	wire        [31:0] w_fld_output_7_dataout_0;
	wire               w_fld_output_7_r_w_0;
	wire               w_fld_output_7_ce_0;
	reg  signed        r_fld_output_7_addr_1;
	reg         [31:0] r_fld_output_7_datain_1;
	wire        [31:0] w_fld_output_7_dataout_1;
	reg                r_fld_output_7_r_w_1;
	wire               w_fld_output_7_ce_1;
	wire signed [ 2:0] w_fld_in_8_addr_0;
	wire        [31:0] w_fld_in_8_datain_0;
	wire        [31:0] w_fld_in_8_dataout_0;
	wire               w_fld_in_8_r_w_0;
	wire               w_fld_in_8_ce_0;
	reg  signed [ 2:0] r_fld_in_8_addr_1;
	reg         [31:0] r_fld_in_8_datain_1;
	wire        [31:0] w_fld_in_8_dataout_1;
	reg                r_fld_in_8_r_w_1;
	wire               w_fld_in_8_ce_1;
	wire signed [ 1:0] w_fld_res_9_addr_0;
	wire        [31:0] w_fld_res_9_datain_0;
	wire        [31:0] w_fld_res_9_dataout_0;
	wire               w_fld_res_9_r_w_0;
	wire               w_fld_res_9_ce_0;
	reg  signed [ 1:0] r_fld_res_9_addr_1;
	reg         [31:0] r_fld_res_9_datain_1;
	wire        [31:0] w_fld_res_9_dataout_1;
	reg                r_fld_res_9_r_w_1;
	wire               w_fld_res_9_ce_1;
	reg         [31:0] r_threadTop_err_10;
	reg         [31:0] r_threadTop_alpha_11;
	reg         [31:0] r_threadTop_sum_12;
	reg         [31:0] r_threadTop_delta_13;
	reg  signed [31:0] r_threadTop_i_14;
	reg  signed [31:0] r_threadTop_j_15;
	reg  signed [31:0] r_threadTop_k_16;
	reg  signed [31:0] r_threadTop_j_17;
	reg  signed [31:0] r_threadTop_k_18;
	reg  signed [31:0] r_threadTop_j_19;
	reg  signed [31:0] r_threadTop_k_20;
	reg  signed [31:0] r_threadTop_j_21;
	reg  signed [31:0] r_threadTop_l_22;
	reg  signed [31:0] r_threadTop_k_23;
	reg  signed [31:0] r_threadTop_j_24;
	reg  signed [31:0] r_threadTop_k_25;
	reg  signed [31:0] r_threadTop_copy0_j_27;
	reg  signed [31:0] r_threadTop_copy0_j_28;
	reg  signed [31:0] r_threadTop_copy0_j_29;
	reg  signed [31:0] r_threadTop_copy0_j_30;
	reg  signed [31:0] r_threadTop_copy1_j_31;
	reg  signed [31:0] r_threadTop_copy0_j_32;
	reg  signed [31:0] r_threadTop_copy1_j_33;
	reg  signed [31:0] r_sys_tmp0_int;
	reg  signed [31:0] r_sys_tmp1_int;
	reg  signed [31:0] r_sys_tmp2_int;
	reg  signed [31:0] r_sys_tmp3_int;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg  signed [31:0] r_sys_tmp4_int;
	reg  signed [31:0] r_sys_tmp5_int;
	reg  signed [31:0] r_sys_tmp6_int;
	reg  signed [31:0] r_sys_tmp7_int;
	reg  signed [31:0] r_sys_tmp8_int;
	reg  signed [31:0] r_sys_tmp9_int;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	wire        [31:0] w_sys_tmp1;
	wire        [31:0] w_sys_tmp3;
	wire signed [31:0] w_sys_tmp7;
	wire signed [31:0] w_sys_tmp10;
	wire signed [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp16;
	wire signed [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp22;
	wire        [31:0] w_sys_tmp35;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp40;
	wire        [31:0] w_sys_tmp43;
	wire        [31:0] w_sys_tmp46;
	wire        [31:0] w_sys_tmp49;
	wire        [31:0] w_sys_tmp52;
	wire        [31:0] w_sys_tmp55;
	wire signed [31:0] w_sys_tmp57;
	wire        [31:0] w_sys_tmp58;
	wire signed [31:0] w_sys_tmp60;
	wire        [31:0] w_sys_tmp61;
	wire        [31:0] w_sys_tmp63;
	wire        [31:0] w_sys_tmp65;
	wire        [31:0] w_sys_tmp68;
	wire        [31:0] w_sys_tmp71;
	wire        [31:0] w_sys_tmp74;
	wire        [31:0] w_sys_tmp75;
	wire               w_sys_tmp76;
	wire signed [31:0] w_sys_tmp77;
	wire               w_sys_tmp79;
	wire        [31:0] w_sys_tmp82;
	wire signed [31:0] w_sys_tmp83;
	wire signed [31:0] w_sys_tmp84;
	wire signed [31:0] w_sys_tmp85;
	wire signed [31:0] w_sys_tmp86;
	wire signed [31:0] w_sys_tmp87;
	wire signed [31:0] w_sys_tmp92;
	wire               w_sys_tmp116;
	wire        [31:0] w_sys_tmp119;
	wire               w_sys_tmp120;
	wire        [31:0] w_sys_tmp123;
	wire        [31:0] w_sys_tmp124;
	wire        [31:0] w_sys_tmp125;
	wire signed [31:0] w_sys_tmp126;
	wire signed [31:0] w_sys_tmp127;
	wire signed [31:0] w_sys_tmp128;
	wire        [31:0] w_sys_tmp129;
	wire signed [31:0] w_sys_tmp130;
	wire signed [31:0] w_sys_tmp131;
	wire        [31:0] w_sys_tmp134;
	wire signed [31:0] w_sys_tmp136;
	wire signed [31:0] w_sys_tmp138;
	wire        [31:0] w_sys_tmp173;
	wire        [31:0] w_sys_tmp174;
	wire        [31:0] w_sys_tmp175;
	wire        [31:0] w_sys_tmp177;
	wire        [31:0] w_sys_tmp178;
	wire        [31:0] w_sys_tmp179;
	wire signed [31:0] w_sys_tmp180;
	wire               w_sys_tmp181;
	wire        [31:0] w_sys_tmp184;
	wire               w_sys_tmp185;
	wire        [31:0] w_sys_tmp188;
	wire        [31:0] w_sys_tmp189;
	wire        [31:0] w_sys_tmp190;
	wire signed [31:0] w_sys_tmp191;
	wire        [31:0] w_sys_tmp192;
	wire signed [31:0] w_sys_tmp193;
	wire signed [31:0] w_sys_tmp194;
	wire        [31:0] w_sys_tmp197;
	wire signed [31:0] w_sys_tmp199;
	wire        [31:0] w_sys_tmp228;
	wire        [31:0] w_sys_tmp229;
	wire        [31:0] w_sys_tmp230;
	wire        [31:0] w_sys_tmp232;
	wire        [31:0] w_sys_tmp233;
	wire        [31:0] w_sys_tmp234;
	wire signed [31:0] w_sys_tmp235;
	wire               w_sys_tmp236;
	wire signed [31:0] w_sys_tmp237;
	wire               w_sys_tmp238;
	wire        [31:0] w_sys_tmp240;
	wire        [31:0] w_sys_tmp241;
	wire        [31:0] w_sys_tmp245;
	wire        [31:0] w_sys_tmp246;
	wire        [31:0] w_sys_tmp247;
	wire signed [31:0] w_sys_tmp248;
	wire        [31:0] w_sys_tmp249;
	wire        [31:0] w_sys_tmp250;
	wire signed [31:0] w_sys_tmp254;
	wire        [31:0] w_sys_tmp255;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp257;
	wire signed [31:0] w_sys_tmp258;
	wire signed [31:0] w_sys_tmp271;
	wire        [31:0] w_sys_tmp273;
	wire signed [31:0] w_sys_tmp274;
	wire               w_sys_tmp335;
	wire signed [31:0] w_sys_tmp336;
	wire        [31:0] w_sys_tmp337;
	wire               w_sys_tmp338;
	wire        [31:0] w_sys_tmp340;
	wire        [31:0] w_sys_tmp341;
	wire signed [31:0] w_sys_tmp344;
	wire        [31:0] w_sys_tmp346;
	wire signed [31:0] w_sys_tmp347;
	wire        [31:0] w_sys_tmp348;
	wire        [31:0] w_sys_tmp349;
	wire signed [31:0] w_sys_tmp351;
	wire               w_sys_tmp352;
	wire        [31:0] w_sys_tmp354;
	wire        [31:0] w_sys_tmp357;
	wire        [31:0] w_sys_tmp358;
	wire        [31:0] w_sys_tmp359;
	wire signed [31:0] w_sys_tmp362;
	wire signed [31:0] w_sys_tmp363;
	wire signed [31:0] w_sys_tmp365;
	wire signed [31:0] w_sys_tmp366;
	wire        [31:0] w_sys_tmp368;
	wire signed [31:0] w_sys_tmp369;
	wire signed [31:0] w_sys_tmp370;
	wire signed [31:0] w_sys_tmp371;
	wire signed [31:0] w_sys_tmp380;
	wire signed [31:0] w_sys_tmp382;
	wire        [31:0] w_sys_tmp384;
	wire signed [31:0] w_sys_tmp385;
	wire signed [31:0] w_sys_tmp387;
	wire        [31:0] w_sys_tmp448;
	wire               w_sys_tmp449;
	wire        [31:0] w_sys_tmp451;
	wire        [31:0] w_sys_tmp452;
	wire        [31:0] w_sys_tmp453;
	wire signed [31:0] w_sys_tmp454;
	wire        [31:0] w_sys_tmp455;
	wire signed [31:0] w_sys_tmp459;
	wire        [31:0] w_sys_tmp460;
	wire        [31:0] w_sys_tmp461;
	wire signed [31:0] w_sys_tmp462;
	wire               w_sys_tmp463;
	wire        [31:0] w_sys_tmp464;
	wire signed [31:0] w_sys_tmp465;
	wire signed [31:0] w_sys_tmp466;
	wire signed [31:0] w_sys_tmp467;
	wire signed [31:0] w_sys_tmp471;
	wire signed [31:0] w_sys_tmp475;
	wire signed [31:0] w_sys_tmp479;
	wire signed [31:0] w_sys_tmp480;
	wire signed [31:0] w_sys_tmp481;
	wire signed [31:0] w_sys_tmp488;
	wire signed [31:0] w_sys_tmp489;
	wire signed [31:0] w_sys_tmp490;
	wire signed [31:0] w_sys_tmp497;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_threadTop_busy = r_sys_threadTop_busy;
	assign w_sys_threadTop_stage_p1 = (r_sys_threadTop_stage + 2'h1);
	assign w_sys_threadTop_step_p1 = (r_sys_threadTop_step + 7'h1);
	assign w_fld_w1_3_addr_0 = 4'sh0;
	assign w_fld_w1_3_datain_0 = 32'h0;
	assign w_fld_w1_3_r_w_0 = 1'h0;
	assign w_fld_w1_3_ce_0 = w_sys_ce;
	assign w_fld_w1_3_ce_1 = w_sys_ce;
	assign w_fld_w2_4_addr_0 = 3'sh0;
	assign w_fld_w2_4_datain_0 = 32'h0;
	assign w_fld_w2_4_r_w_0 = 1'h0;
	assign w_fld_w2_4_ce_0 = w_sys_ce;
	assign w_fld_w2_4_ce_1 = w_sys_ce;
	assign w_fld_input_5_addr_0 = 1'sh0;
	assign w_fld_input_5_datain_0 = 32'h0;
	assign w_fld_input_5_r_w_0 = 1'h0;
	assign w_fld_input_5_ce_0 = w_sys_ce;
	assign w_fld_input_5_ce_1 = w_sys_ce;
	assign w_fld_hidden_6_addr_0 = 3'sh0;
	assign w_fld_hidden_6_datain_0 = 32'h0;
	assign w_fld_hidden_6_r_w_0 = 1'h0;
	assign w_fld_hidden_6_ce_0 = w_sys_ce;
	assign w_fld_hidden_6_ce_1 = w_sys_ce;
	assign w_fld_output_7_addr_0 = 1'sh0;
	assign w_fld_output_7_datain_0 = 32'h0;
	assign w_fld_output_7_r_w_0 = 1'h0;
	assign w_fld_output_7_ce_0 = w_sys_ce;
	assign w_fld_output_7_ce_1 = w_sys_ce;
	assign w_fld_in_8_addr_0 = 3'sh0;
	assign w_fld_in_8_datain_0 = 32'h0;
	assign w_fld_in_8_r_w_0 = 1'h0;
	assign w_fld_in_8_ce_0 = w_sys_ce;
	assign w_fld_in_8_ce_1 = w_sys_ce;
	assign w_fld_res_9_addr_0 = 2'sh0;
	assign w_fld_res_9_datain_0 = 32'h0;
	assign w_fld_res_9_r_w_0 = 1'h0;
	assign w_fld_res_9_ce_0 = w_sys_ce;
	assign w_fld_res_9_ce_1 = w_sys_ce;
	assign w_sys_tmp1 = 32'h0;
	assign w_sys_tmp3 = 32'h3f800000;
	assign w_sys_tmp7 = 32'sh00000002;
	assign w_sys_tmp10 = 32'sh00000003;
	assign w_sys_tmp13 = 32'sh00000004;
	assign w_sys_tmp16 = 32'sh00000005;
	assign w_sys_tmp19 = 32'sh00000006;
	assign w_sys_tmp22 = 32'sh00000007;
	assign w_sys_tmp35 = 32'hbc0c825a;
	assign w_sys_tmp37 = 32'h3d4d320d;
	assign w_sys_tmp40 = 32'hbd4d74b0;
	assign w_sys_tmp43 = 32'hbdc24c38;
	assign w_sys_tmp46 = 32'h3d4b55a3;
	assign w_sys_tmp49 = 32'hbd9d6bc6;
	assign w_sys_tmp52 = 32'hbd0b991f;
	assign w_sys_tmp55 = 32'h3d5b1cfd;
	assign w_sys_tmp57 = 32'sh00000008;
	assign w_sys_tmp58 = 32'h3dc048ab;
	assign w_sys_tmp60 = 32'sh00000009;
	assign w_sys_tmp61 = 32'hbb6d0bb3;
	assign w_sys_tmp63 = 32'h3bc88e80;
	assign w_sys_tmp65 = 32'hbda4d7e7;
	assign w_sys_tmp68 = 32'h3cda20ed;
	assign w_sys_tmp71 = 32'hbc6f47b3;
	assign w_sys_tmp74 = 32'hbd625c80;
	assign w_sys_tmp75 = 32'h3dcccccd;
	assign w_sys_tmp76 = (r_threadTop_i_14 < w_sys_tmp77);
	assign w_sys_tmp77 = 32'sh00000004;
	assign w_sys_tmp79 = (r_threadTop_j_15 < r_fld_N_INPUT_0);
	assign w_sys_tmp82 = w_fld_in_8_dataout_1;
	assign w_sys_tmp83 = (w_sys_tmp84 + r_threadTop_copy0_j_27);
	assign w_sys_tmp84 = (w_sys_tmp85 * r_threadTop_i_14);
	assign w_sys_tmp85 = 32'sh00000002;
	assign w_sys_tmp86 = (r_threadTop_copy0_j_27 + w_sys_intOne);
	assign w_sys_tmp87 = (r_threadTop_j_15 + w_sys_intOne);
	assign w_sys_tmp92 = w_sys_tmp86;
	assign w_sys_tmp116 = (r_threadTop_k_16 < r_fld_N_HIDDEN_1);
	assign w_sys_tmp119 = 32'h0;
	assign w_sys_tmp120 = (r_threadTop_j_17 < r_fld_N_INPUT_0);
	assign w_sys_tmp123 = w_ip_AddFloat_result_0;
	assign w_sys_tmp124 = w_ip_MultFloat_product_0;
	assign w_sys_tmp125 = w_fld_w1_3_dataout_1;
	assign w_sys_tmp126 = (w_sys_tmp127 + r_threadTop_k_16);
	assign w_sys_tmp127 = (w_sys_tmp128 * r_threadTop_j_17);
	assign w_sys_tmp128 = 32'sh00000005;
	assign w_sys_tmp129 = w_fld_input_5_dataout_1;
	assign w_sys_tmp130 = (r_threadTop_copy0_j_28 + w_sys_intOne);
	assign w_sys_tmp131 = (r_threadTop_j_17 + w_sys_intOne);
	assign w_sys_tmp134 = w_fld_hidden_6_dataout_1;
	assign w_sys_tmp136 = (w_sys_tmp128 * w_sys_tmp138);
	assign w_sys_tmp138 = w_sys_tmp131;
	assign w_sys_tmp173 = w_ip_DivFloat_quotient_0;
	assign w_sys_tmp174 = 32'h3f800000;
	assign w_sys_tmp175 = w_ip_AddFloat_result_0;
	assign w_sys_tmp177 = w_ip_exp_result_0;
	assign w_sys_tmp178 = ( -w_sys_tmp179 );
	assign w_sys_tmp179 = w_fld_hidden_6_dataout_1;
	assign w_sys_tmp180 = (r_threadTop_k_16 + w_sys_intOne);
	assign w_sys_tmp181 = (r_threadTop_k_18 < r_fld_N_OUTPUT_2);
	assign w_sys_tmp184 = 32'h0;
	assign w_sys_tmp185 = (r_threadTop_j_19 < r_fld_N_HIDDEN_1);
	assign w_sys_tmp188 = w_ip_AddFloat_result_0;
	assign w_sys_tmp189 = w_ip_MultFloat_product_0;
	assign w_sys_tmp190 = w_fld_w2_4_dataout_1;
	assign w_sys_tmp191 = (r_threadTop_j_19 + r_threadTop_k_18);
	assign w_sys_tmp192 = w_fld_hidden_6_dataout_1;
	assign w_sys_tmp193 = (r_threadTop_copy0_j_29 + w_sys_intOne);
	assign w_sys_tmp194 = (r_threadTop_j_19 + w_sys_intOne);
	assign w_sys_tmp197 = w_fld_output_7_dataout_1;
	assign w_sys_tmp199 = w_sys_tmp194;
	assign w_sys_tmp228 = w_ip_DivFloat_quotient_0;
	assign w_sys_tmp229 = 32'h3f800000;
	assign w_sys_tmp230 = w_ip_AddFloat_result_0;
	assign w_sys_tmp232 = w_ip_exp_result_1;
	assign w_sys_tmp233 = ( -w_sys_tmp234 );
	assign w_sys_tmp234 = w_fld_output_7_dataout_1;
	assign w_sys_tmp235 = (r_threadTop_k_18 + w_sys_intOne);
	assign w_sys_tmp236 = (r_threadTop_k_20 < r_fld_N_OUTPUT_2);
	assign w_sys_tmp237 = (r_threadTop_k_20 + w_sys_intOne);
	assign w_sys_tmp238 = (r_threadTop_j_21 < r_fld_N_HIDDEN_1);
	assign w_sys_tmp240 = w_ip_MultFloat_product_0;
	assign w_sys_tmp241 = ( -r_threadTop_alpha_11 );
	assign w_sys_tmp245 = ( -w_sys_tmp246 );
	assign w_sys_tmp246 = w_ip_AddFloat_result_0;
	assign w_sys_tmp247 = w_fld_res_9_dataout_1;
	assign w_sys_tmp248 = (r_threadTop_i_14 + r_threadTop_k_20);
	assign w_sys_tmp249 = w_fld_output_7_dataout_1;
	assign w_sys_tmp250 = 32'h3f800000;
	assign w_sys_tmp254 = (r_threadTop_copy0_j_30 + r_threadTop_k_20);
	assign w_sys_tmp255 = w_sys_tmp240;
	assign w_sys_tmp256 = (r_threadTop_copy0_j_30 + w_sys_intOne);
	assign w_sys_tmp257 = (r_threadTop_copy1_j_31 + w_sys_intOne);
	assign w_sys_tmp258 = (r_threadTop_j_21 + w_sys_intOne);
	assign w_sys_tmp271 = w_sys_tmp257;
	assign w_sys_tmp273 = w_fld_w2_4_dataout_1;
	assign w_sys_tmp274 = w_sys_tmp256;
	assign w_sys_tmp335 = (r_threadTop_l_22 < r_fld_N_HIDDEN_1);
	assign w_sys_tmp336 = (r_threadTop_l_22 + w_sys_intOne);
	assign w_sys_tmp337 = 32'h0;
	assign w_sys_tmp338 = (r_threadTop_k_23 < r_fld_N_OUTPUT_2);
	assign w_sys_tmp340 = w_ip_AddFloat_result_0;
	assign w_sys_tmp341 = w_ip_MultFloat_product_0;
	assign w_sys_tmp344 = (r_threadTop_l_22 + r_threadTop_k_23);
	assign w_sys_tmp346 = w_fld_res_9_dataout_1;
	assign w_sys_tmp347 = (r_threadTop_i_14 + r_threadTop_k_23);
	assign w_sys_tmp348 = w_fld_output_7_dataout_1;
	assign w_sys_tmp349 = 32'h3f800000;
	assign w_sys_tmp351 = (r_threadTop_k_23 + w_sys_intOne);
	assign w_sys_tmp352 = (r_threadTop_j_24 < r_fld_N_INPUT_0);
	assign w_sys_tmp354 = w_ip_MultFloat_product_0;
	assign w_sys_tmp357 = w_fld_hidden_6_dataout_1;
	assign w_sys_tmp358 = w_ip_AddFloat_result_0;
	assign w_sys_tmp359 = 32'h3f800000;
	assign w_sys_tmp362 = (w_sys_tmp363 * r_threadTop_copy1_j_33);
	assign w_sys_tmp363 = 32'sh00000005;
	assign w_sys_tmp365 = (w_sys_tmp366 + r_threadTop_l_22);
	assign w_sys_tmp366 = (w_sys_tmp363 * r_threadTop_copy0_j_32);
	assign w_sys_tmp368 = w_sys_tmp354;
	assign w_sys_tmp369 = (r_threadTop_copy0_j_32 + w_sys_intOne);
	assign w_sys_tmp370 = (r_threadTop_copy1_j_33 + w_sys_intOne);
	assign w_sys_tmp371 = (r_threadTop_j_24 + w_sys_intOne);
	assign w_sys_tmp380 = (w_sys_tmp363 * w_sys_tmp382);
	assign w_sys_tmp382 = w_sys_tmp370;
	assign w_sys_tmp384 = w_fld_w1_3_dataout_1;
	assign w_sys_tmp385 = (w_sys_tmp363 * w_sys_tmp387);
	assign w_sys_tmp387 = w_sys_tmp369;
	assign w_sys_tmp448 = 32'h0;
	assign w_sys_tmp449 = (r_threadTop_k_25 < r_fld_N_OUTPUT_2);
	assign w_sys_tmp451 = w_ip_AddFloat_result_0;
	assign w_sys_tmp452 = w_ip_MultFloat_product_0;
	assign w_sys_tmp453 = w_fld_res_9_dataout_1;
	assign w_sys_tmp454 = (r_threadTop_i_14 + r_threadTop_k_25);
	assign w_sys_tmp455 = w_fld_output_7_dataout_1;
	assign w_sys_tmp459 = (r_threadTop_k_25 + w_sys_intOne);
	assign w_sys_tmp460 = w_ip_MultFloat_product_0;
	assign w_sys_tmp461 = 32'h3f000000;
	assign w_sys_tmp462 = (r_threadTop_i_14 + w_sys_intOne);
	assign w_sys_tmp463 = w_ip_CompareFloatLT_result_0;
	assign w_sys_tmp464 = 32'h3a83126f;
	assign w_sys_tmp465 = 32'sh00000002;
	assign w_sys_tmp466 = 32'sh00000005;
	assign w_sys_tmp467 = (w_sys_tmp84 + w_sys_tmp92);
	assign w_sys_tmp471 = (w_sys_tmp136 + r_threadTop_k_16);
	assign w_sys_tmp475 = (w_sys_tmp199 + r_threadTop_k_18);
	assign w_sys_tmp479 = (r_threadTop_copy1_j_31 + r_threadTop_k_20);
	assign w_sys_tmp480 = (w_sys_tmp271 + r_threadTop_k_20);
	assign w_sys_tmp481 = (w_sys_tmp274 + r_threadTop_k_20);
	assign w_sys_tmp488 = (w_sys_tmp362 + r_threadTop_l_22);
	assign w_sys_tmp489 = (w_sys_tmp380 + r_threadTop_l_22);
	assign w_sys_tmp490 = (w_sys_tmp385 + r_threadTop_l_22);
	assign w_sys_tmp497 = (r_threadTop_i_14 + r_threadTop_k_25);


	DualPortRAM #(.DWIDTH(32), .AWIDTH(4), .WORDS(10) )
		dpram_w1_3(
			.clk (clock),
			.ce_0 (w_fld_w1_3_ce_0),
			.addr_0 (w_fld_w1_3_addr_0),
			.datain_0 (w_fld_w1_3_datain_0),
			.dataout_0 (w_fld_w1_3_dataout_0),
			.r_w_0 (w_fld_w1_3_r_w_0),
			.ce_1 (w_fld_w1_3_ce_1),
			.addr_1 (r_fld_w1_3_addr_1),
			.datain_1 (r_fld_w1_3_datain_1),
			.dataout_1 (w_fld_w1_3_dataout_1),
			.r_w_1 (r_fld_w1_3_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(3), .WORDS(5) )
		dpram_w2_4(
			.clk (clock),
			.ce_0 (w_fld_w2_4_ce_0),
			.addr_0 (w_fld_w2_4_addr_0),
			.datain_0 (w_fld_w2_4_datain_0),
			.dataout_0 (w_fld_w2_4_dataout_0),
			.r_w_0 (w_fld_w2_4_r_w_0),
			.ce_1 (w_fld_w2_4_ce_1),
			.addr_1 (r_fld_w2_4_addr_1),
			.datain_1 (r_fld_w2_4_datain_1),
			.dataout_1 (w_fld_w2_4_dataout_1),
			.r_w_1 (r_fld_w2_4_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(1), .WORDS(2) )
		dpram_input_5(
			.clk (clock),
			.ce_0 (w_fld_input_5_ce_0),
			.addr_0 (w_fld_input_5_addr_0),
			.datain_0 (w_fld_input_5_datain_0),
			.dataout_0 (w_fld_input_5_dataout_0),
			.r_w_0 (w_fld_input_5_r_w_0),
			.ce_1 (w_fld_input_5_ce_1),
			.addr_1 (r_fld_input_5_addr_1),
			.datain_1 (r_fld_input_5_datain_1),
			.dataout_1 (w_fld_input_5_dataout_1),
			.r_w_1 (r_fld_input_5_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(3), .WORDS(5) )
		dpram_hidden_6(
			.clk (clock),
			.ce_0 (w_fld_hidden_6_ce_0),
			.addr_0 (w_fld_hidden_6_addr_0),
			.datain_0 (w_fld_hidden_6_datain_0),
			.dataout_0 (w_fld_hidden_6_dataout_0),
			.r_w_0 (w_fld_hidden_6_r_w_0),
			.ce_1 (w_fld_hidden_6_ce_1),
			.addr_1 (r_fld_hidden_6_addr_1),
			.datain_1 (r_fld_hidden_6_datain_1),
			.dataout_1 (w_fld_hidden_6_dataout_1),
			.r_w_1 (r_fld_hidden_6_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(1), .WORDS(1) )
		dpram_output_7(
			.clk (clock),
			.ce_0 (w_fld_output_7_ce_0),
			.addr_0 (w_fld_output_7_addr_0),
			.datain_0 (w_fld_output_7_datain_0),
			.dataout_0 (w_fld_output_7_dataout_0),
			.r_w_0 (w_fld_output_7_r_w_0),
			.ce_1 (w_fld_output_7_ce_1),
			.addr_1 (r_fld_output_7_addr_1),
			.datain_1 (r_fld_output_7_datain_1),
			.dataout_1 (w_fld_output_7_dataout_1),
			.r_w_1 (r_fld_output_7_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(3), .WORDS(8) )
		dpram_in_8(
			.clk (clock),
			.ce_0 (w_fld_in_8_ce_0),
			.addr_0 (w_fld_in_8_addr_0),
			.datain_0 (w_fld_in_8_datain_0),
			.dataout_0 (w_fld_in_8_dataout_0),
			.r_w_0 (w_fld_in_8_r_w_0),
			.ce_1 (w_fld_in_8_ce_1),
			.addr_1 (r_fld_in_8_addr_1),
			.datain_1 (r_fld_in_8_datain_1),
			.dataout_1 (w_fld_in_8_dataout_1),
			.r_w_1 (r_fld_in_8_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(2), .WORDS(4) )
		dpram_res_9(
			.clk (clock),
			.ce_0 (w_fld_res_9_ce_0),
			.addr_0 (w_fld_res_9_addr_0),
			.datain_0 (w_fld_res_9_datain_0),
			.dataout_0 (w_fld_res_9_dataout_0),
			.r_w_0 (w_fld_res_9_r_w_0),
			.ce_1 (w_fld_res_9_ce_1),
			.addr_1 (r_fld_res_9_addr_1),
			.datain_1 (r_fld_res_9_datain_1),
			.dataout_1 (w_fld_res_9_dataout_1),
			.r_w_1 (r_fld_res_9_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	DivFloat
		DivFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_DivFloat_dividend_0),
			.b (r_ip_DivFloat_divisor_0),
			.result (w_ip_DivFloat_quotient_0)
		);

	CompareFloatLT
		CompareFloatLT_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_CompareFloatLT_portA_0),
			.b (r_ip_CompareFloatLT_portB_0),
			.result (w_ip_CompareFloatLT_result_0)
		);

	exp
		exp_inst_0(
			.clk (clock),
			.nD (r_ip_exp_newData_0),
			.i (r_ip_exp_i_0),	// in 32bit
			.out (w_ip_exp_result_0)	// out 32bit
		);

	exp
		exp_inst_1(
			.clk (clock),
			.nD (r_ip_exp_newData_1),
			.i (r_ip_exp_i_1),	// in 32bit
			.out (w_ip_exp_result_1)	// out 32bit
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hf) || (r_sys_threadTop_step==7'h17) || (r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h27)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp134;

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp3_float;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp174;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_threadTop_step==7'hf) || (r_sys_threadTop_step==7'h17) || (r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h27)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp197;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp229;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h23) || (r_sys_threadTop_step==7'h2b) || (r_sys_threadTop_step==7'h33) || (r_sys_threadTop_step==7'h3b)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp273;

									end
									else
									if((r_sys_threadTop_step==7'he)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp247;

									end
									else
									if((r_sys_threadTop_step==7'h5) || (r_sys_threadTop_step==7'hb)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_threadTop_step==7'h4) || (r_sys_threadTop_step==7'h7) || (r_sys_threadTop_step==7'ha) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h10)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp250;

									end
									else
									if((r_sys_threadTop_step==7'h1b)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp6_float;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h4)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp349;

									end
									else
									if((r_sys_threadTop_step==7'h16)) begin
										r_ip_AddFloat_portA_0 <= r_threadTop_sum_12;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp346;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h27) || (r_sys_threadTop_step==7'h2f) || (r_sys_threadTop_step==7'h37)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp384;

									end
									else
									if((r_sys_threadTop_step==7'h17)) begin
										r_ip_AddFloat_portA_0 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_threadTop_step==7'h3) || (r_sys_threadTop_step==7'h5) || (r_sys_threadTop_step==7'h7) || (r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hb)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp359;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hd)) begin
										r_ip_AddFloat_portA_0 <= r_threadTop_err_10;

									end
									else
									if((r_sys_threadTop_step==7'h2) || (r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp453;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hf)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp124;

									end
									else
									if((r_sys_threadTop_step==7'h1f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_threadTop_step==7'h27)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_threadTop_step==7'h17)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp177;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hf)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'h1f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_threadTop_step==7'h27)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp189;

									end
									else
									if((r_sys_threadTop_step==7'h17)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp232;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp249[31], w_sys_tmp249[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'hb)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp249[31], w_sys_tmp249[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp249[31], w_sys_tmp249[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h5)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp249[31], w_sys_tmp249[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp249[31], w_sys_tmp249[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp249[31], w_sys_tmp249[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp249[31], w_sys_tmp249[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp249[31], w_sys_tmp249[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h23) || (r_sys_threadTop_step==7'h33)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_threadTop_step==7'ha)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp249[31], w_sys_tmp249[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h3b)) begin
										r_ip_AddFloat_portB_0 <= r_threadTop_delta_13;

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp249[31], w_sys_tmp249[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h2b)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_threadTop_step==7'h1b)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp255;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp348[31], w_sys_tmp348[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp348[31], w_sys_tmp348[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h16)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp341;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp357[31], w_sys_tmp357[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h5)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp357[31], w_sys_tmp357[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'hb)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp357[31], w_sys_tmp357[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp357[31], w_sys_tmp357[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h2f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'h17)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp368;

									end
									else
									if((r_sys_threadTop_step==7'h9)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp357[31], w_sys_tmp357[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'h27)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_threadTop_step==7'h37)) begin
										r_ip_AddFloat_portB_0 <= r_threadTop_delta_13;

									end
									else
									if((r_sys_threadTop_step==7'h1f)) begin
										r_ip_AddFloat_portB_0 <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp455[31], w_sys_tmp455[30:0] };

									end
									else
									if((r_sys_threadTop_step==7'hd)) begin
										r_ip_AddFloat_portB_0 <= w_sys_tmp452;

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp455[31], w_sys_tmp455[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp125;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp190;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7) || (r_sys_threadTop_step==7'ha) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h10) || (r_sys_threadTop_step==7'h13)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp245;

									end
									else
									if((r_sys_threadTop_step==7'h16) || (r_sys_threadTop_step==7'h19) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h22)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp241;

									end
									else
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'hf) || (r_sys_threadTop_step==7'h11) || (r_sys_threadTop_step==7'h12) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h17) || (r_sys_threadTop_step==7'h18) || (r_sys_threadTop_step==7'h1a) || (r_sys_threadTop_step==7'h1d)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp240;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'h11)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp341;

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'hd<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h16) || (r_sys_threadTop_step==7'h18) || (r_sys_threadTop_step==7'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp354;

									end
									else
									if((r_sys_threadTop_step==7'h8) || (r_sys_threadTop_step==7'ha) || (r_sys_threadTop_step==7'hc)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'h2) || (r_sys_threadTop_step==7'h4) || (r_sys_threadTop_step==7'h6) || (r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hb)) begin
										r_ip_MultFloat_multiplicand_0 <= r_threadTop_alpha_11;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp6_float;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_ip_MultFloat_multiplicand_0 <= r_threadTop_err_10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp129;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp192;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'ha) || (r_sys_threadTop_step==7'h10)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_threadTop_step==7'h16) || (r_sys_threadTop_step==7'h19) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h1f) || (r_sys_threadTop_step==7'h22)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp240;

									end
									else
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'hf) || (r_sys_threadTop_step==7'h12) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h18)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_threadTop_step==7'h11)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_threadTop_step==7'h17)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_threadTop_step==7'h14)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_threadTop_step==7'h1d)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_threadTop_step==7'h7) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h13)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp9_float;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp340;

									end
									else
									if((r_sys_threadTop_step==7'h11)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_threadTop_step==7'hc)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2) || (r_sys_threadTop_step==7'h4) || (r_sys_threadTop_step==7'h6)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp357;

									end
									else
									if((r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hb)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_threadTop_step==7'hd)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_threadTop_step==7'h12) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h16) || (r_sys_threadTop_step==7'h18) || (r_sys_threadTop_step==7'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_threadTop_sum_12;

									end
									else
									if((r_sys_threadTop_step==7'h15)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_threadTop_step==7'h8) || (r_sys_threadTop_step==7'ha) || (r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'he) || (r_sys_threadTop_step==7'h10)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp358;

									end
									else
									if((r_sys_threadTop_step==7'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_threadTop_step==7'h13)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_threadTop_step==7'h11)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp6_float;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp451;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp461;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_DivFloat_dividend_0 <= w_sys_tmp174;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_DivFloat_dividend_0 <= w_sys_tmp229;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_DivFloat_divisor_0 <= w_sys_tmp175;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_ip_DivFloat_divisor_0 <= w_sys_tmp230;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h51: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_ip_CompareFloatLT_portA_0 <= r_threadTop_err_10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h51: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_ip_CompareFloatLT_portB_0 <= w_sys_tmp464;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_exp_i_0 <= w_sys_tmp178;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_exp_newData_0 <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_exp_i_1 <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_ip_exp_newData_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_threadTop_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h55: begin
							r_sys_processing_methodID <= r_sys_threadTop_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h0: begin
							r_sys_threadTop_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h9)) begin
										r_sys_threadTop_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_boolFalse) ? 7'h7 : 7'h55);

									end
								end

							endcase
						end

						7'h7: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h8;

									end
								end

							endcase
						end

						7'h8: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp76) ? 7'hc : 7'h51);

									end
								end

							endcase
						end

						7'hc: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'hd;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp79) ? 7'h10 : 7'h12);

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_threadTop_phase <= 7'hd;

									end
								end

							endcase
						end

						7'h12: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h13;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp116) ? 7'h16 : 7'h1f);

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h18;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h19;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp120) ? 7'h1c : 7'h1d);

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_phase <= 7'h19;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_phase <= 7'h13;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h20;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp181) ? 7'h23 : 7'h2c);

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h25;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h26;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp185) ? 7'h29 : 7'h2a);

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_phase <= 7'h26;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_phase <= 7'h20;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp236) ? 7'h31 : 7'h37);

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h32;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp238) ? 7'h35 : 7'h2e);

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h40)) begin
										r_sys_threadTop_phase <= 7'h32;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h38;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp335) ? 7'h3b : 7'h48);

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h38;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h3d;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h3e;

									end
								end

							endcase
						end

						7'h3e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp338) ? 7'h41 : 7'h43);

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b)) begin
										r_sys_threadTop_phase <= 7'h3e;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h44;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp352) ? 7'h47 : 7'h39);

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3c)) begin
										r_sys_threadTop_phase <= 7'h44;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h4a;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= 7'h4b;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp449) ? 7'h4e : 7'h4f);

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h12)) begin
										r_sys_threadTop_phase <= 7'h4b;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_sys_threadTop_phase <= 7'h8;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_threadTop_phase <= ((w_sys_tmp463) ? 7'h53 : 7'h4);

									end
								end

							endcase
						end

						7'h53: begin
							r_sys_threadTop_phase <= 7'h55;
						end

						7'h55: begin
							r_sys_threadTop_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_stage <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h9)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h7: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h8: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'hc: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h12: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h40)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h3e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= w_sys_threadTop_stage_p1;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3c)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h12)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_threadTop_stage <= 2'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h9)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h8)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h7: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h8: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'hc: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h5)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h12: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h2b)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h25)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h1f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h25: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2c)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h2b)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h25)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h31: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h40)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3f)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h37: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h1a)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h43: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h44: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3c)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3b)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_threadTop_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h12)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h11)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

						7'h51: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_threadTop_step <= 7'h0;

									end
									else
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1) || (r_sys_threadTop_step==7'h2)) begin
										r_sys_threadTop_step <= w_sys_threadTop_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_threadTop_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_threadTop_busy <= ((i_threadTop_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h0: begin
							r_sys_threadTop_busy <= w_sys_boolTrue;
						end

						7'h55: begin
							r_sys_threadTop_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_N_INPUT_0 <= w_sys_tmp465;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_N_HIDDEN_1 <= w_sys_tmp466;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_N_OUTPUT_2 <= w_sys_intOne;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_w1_3_addr_1 <= 4'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp16[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_intZero[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h8)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp57[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp7[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_intOne[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h9)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp60[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp22[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp13[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp10[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h6)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp19[3:0] );

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp126[3:0] );

									end
									else
									if((7'h1<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_w1_3_addr_1 <= $signed( r_sys_tmp1_int[3:0] );

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1d)) begin
										r_fld_w1_3_addr_1 <= $signed( r_sys_tmp2_int[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h25)) begin
										r_fld_w1_3_addr_1 <= $signed( r_sys_tmp5_int[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w1_3_addr_1 <= $signed( w_sys_tmp365[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h34)) begin
										r_fld_w1_3_addr_1 <= $signed( r_sys_tmp4_int[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h24)) begin
										r_fld_w1_3_addr_1 <= $signed( r_sys_tmp1_int[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h3c)) begin
										r_fld_w1_3_addr_1 <= $signed( r_sys_tmp7_int[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h1c)) begin
										r_fld_w1_3_addr_1 <= $signed( r_sys_tmp0_int[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h35)) begin
										r_fld_w1_3_addr_1 <= $signed( r_sys_tmp6_int[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h2c)) begin
										r_fld_w1_3_addr_1 <= $signed( r_sys_tmp9_int[3:0] );

									end
									else
									if((r_sys_threadTop_step==7'h2d)) begin
										r_fld_w1_3_addr_1 <= $signed( r_sys_tmp8_int[3:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp35;

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp46;

									end
									else
									if((r_sys_threadTop_step==7'h8)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp58;

									end
									else
									if((r_sys_threadTop_step==7'h9)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp61;

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp55;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp40;

									end
									else
									if((r_sys_threadTop_step==7'h5)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp49;

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp43;

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp37;

									end
									else
									if((r_sys_threadTop_step==7'h6)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp52;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c) || (r_sys_threadTop_step==7'h34) || (r_sys_threadTop_step==7'h3c)) begin
										r_fld_w1_3_datain_1 <= w_sys_tmp358;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_w1_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h9)) begin
										r_fld_w1_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_w1_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h25) || (r_sys_threadTop_step==7'h2d) || (r_sys_threadTop_step==7'h35)) begin
										r_fld_w1_3_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c) || (r_sys_threadTop_step==7'h34) || (r_sys_threadTop_step==7'h3c)) begin
										r_fld_w1_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h55: begin
							r_fld_w1_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_w2_4_addr_1 <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_intZero[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp7[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_intOne[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp13[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp10[2:0] );

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h1<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_w2_4_addr_1 <= $signed( r_sys_tmp3_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp191[2:0] );

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h31)) begin
										r_fld_w2_4_addr_1 <= $signed( r_sys_tmp2_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h38)) begin
										r_fld_w2_4_addr_1 <= $signed( r_sys_tmp3_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h30)) begin
										r_fld_w2_4_addr_1 <= $signed( r_sys_tmp5_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp254[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h29)) begin
										r_fld_w2_4_addr_1 <= $signed( r_sys_tmp4_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h40)) begin
										r_fld_w2_4_addr_1 <= $signed( r_sys_tmp1_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h28)) begin
										r_fld_w2_4_addr_1 <= $signed( r_sys_tmp7_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h39)) begin
										r_fld_w2_4_addr_1 <= $signed( r_sys_tmp0_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h20)) begin
										r_fld_w2_4_addr_1 <= $signed( r_sys_tmp6_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h21)) begin
										r_fld_w2_4_addr_1 <= $signed( r_sys_tmp8_int[2:0] );

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w2_4_addr_1 <= $signed( w_sys_tmp344[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_fld_w2_4_datain_1 <= w_sys_tmp71;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_fld_w2_4_datain_1 <= w_sys_tmp68;

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w2_4_datain_1 <= w_sys_tmp63;

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_fld_w2_4_datain_1 <= w_sys_tmp74;

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_w2_4_datain_1 <= w_sys_tmp65;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h20) || (r_sys_threadTop_step==7'h28) || (r_sys_threadTop_step==7'h30) || (r_sys_threadTop_step==7'h38) || (r_sys_threadTop_step==7'h40)) begin
										r_fld_w2_4_datain_1 <= w_sys_tmp246;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_w2_4_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_w2_4_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_w2_4_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h21) || (r_sys_threadTop_step==7'h29) || (r_sys_threadTop_step==7'h31) || (r_sys_threadTop_step==7'h39)) begin
										r_fld_w2_4_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTop_step==7'h20) || (r_sys_threadTop_step==7'h28) || (r_sys_threadTop_step==7'h30) || (r_sys_threadTop_step==7'h38) || (r_sys_threadTop_step==7'h40)) begin
										r_fld_w2_4_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_w2_4_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h55: begin
							r_fld_w2_4_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_input_5_addr_1 <= 1'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3) || (r_sys_threadTop_step==7'h6)) begin
										r_fld_input_5_addr_1 <= $signed( r_sys_tmp2_int[0:0] );

									end
									else
									if((r_sys_threadTop_step==7'h2) || (r_sys_threadTop_step==7'h5)) begin
										r_fld_input_5_addr_1 <= $signed( r_sys_tmp1_int[0:0] );

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_fld_input_5_addr_1 <= $signed( r_sys_tmp0_int[0:0] );

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_input_5_addr_1 <= $signed( r_threadTop_copy0_j_28[0:0] );

									end
									else
									if((7'h1<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_input_5_addr_1 <= $signed( r_sys_tmp0_int[0:0] );

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h1<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_input_5_addr_1 <= $signed( r_sys_tmp3_int[0:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_input_5_addr_1 <= $signed( r_threadTop_j_24[0:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_fld_input_5_datain_1 <= w_sys_tmp82;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_input_5_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h2<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h6)) begin
										r_fld_input_5_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_input_5_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_input_5_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h55: begin
							r_fld_input_5_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_hidden_6_addr_1 <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h16: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_k_16[2:0] );

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h25) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_k_16[2:0] );

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_sys_tmp2_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_i_14[2:0] );

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h1<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_sys_tmp2_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_copy0_j_29[2:0] );

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_j_21[2:0] );

									end
									else
									if((7'h1<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_sys_tmp9_int[2:0] );

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h9)) begin
										r_fld_hidden_6_addr_1 <= $signed( r_threadTop_l_22[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h16: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_datain_1 <= w_sys_tmp119;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_hidden_6_datain_1 <= w_sys_tmp123;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_hidden_6_datain_1 <= w_sys_tmp173;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h16: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h25)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h9)) begin
										r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h55: begin
							r_fld_hidden_6_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_output_7_addr_1 <= 1'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_18[0:0] );

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h25) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_18[0:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_output_7_addr_1 <= $signed( r_sys_tmp0_int[0:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_18[0:0] );

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'he)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_20[0:0] );

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_output_7_addr_1 <= $signed( r_sys_tmp5_int[0:0] );

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_fld_output_7_addr_1 <= $signed( r_sys_tmp4_int[0:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_23[0:0] );

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_addr_1 <= $signed( r_threadTop_k_25[0:0] );

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_output_7_addr_1 <= $signed( r_sys_tmp6_int[0:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_datain_1 <= w_sys_tmp184;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_output_7_datain_1 <= w_sys_tmp188;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_output_7_datain_1 <= w_sys_tmp228;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_output_7_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h23: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'hd) || (r_sys_threadTop_step==7'h15) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h25)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'h14) || (r_sys_threadTop_step==7'h1c) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h2c)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_threadTop_step==7'h26)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'he)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1) || (r_sys_threadTop_step==7'h2)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1)) begin
										r_fld_output_7_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h55: begin
							r_fld_output_7_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_in_8_addr_1 <= 3'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp16[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_intZero[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp7[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_intOne[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h7)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp22[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp13[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp10[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h6)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp19[2:0] );

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h1<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_in_8_addr_1 <= $signed( r_sys_tmp3_int[2:0] );

									end
									else
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_in_8_addr_1 <= $signed( w_sys_tmp83[2:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1) || (r_sys_threadTop_step==7'h2) || (r_sys_threadTop_step==7'h5)) begin
										r_fld_in_8_datain_1 <= w_sys_tmp3;

									end
									else
									if((r_sys_threadTop_step==7'h3) || (r_sys_threadTop_step==7'h4) || (r_sys_threadTop_step==7'h6) || (r_sys_threadTop_step==7'h7)) begin
										r_fld_in_8_datain_1 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_in_8_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h7)) begin
										r_fld_in_8_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_in_8_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h55: begin
							r_fld_in_8_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_res_9_addr_1 <= 2'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_intZero[1:0] );

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_tmp7[1:0] );

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_intOne[1:0] );

									end
									else
									if((r_sys_threadTop_step==7'h3)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_tmp10[1:0] );

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_tmp248[1:0] );

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_tmp347[1:0] );

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_res_9_addr_1 <= $signed( w_sys_tmp454[1:0] );

									end
									else
									if((r_sys_threadTop_step==7'h1)) begin
										r_fld_res_9_addr_1 <= $signed( r_sys_tmp7_int[1:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1) || (r_sys_threadTop_step==7'h2)) begin
										r_fld_res_9_datain_1 <= w_sys_tmp3;

									end
									else
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h3)) begin
										r_fld_res_9_datain_1 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_res_9_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3)) begin
										r_fld_res_9_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_fld_res_9_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_fld_res_9_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h1)) begin
										r_fld_res_9_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h55: begin
							r_fld_res_9_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_err_10 <= w_sys_tmp1;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_err_10 <= w_sys_tmp448;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h12)) begin
										r_threadTop_err_10 <= w_sys_tmp451;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_threadTop_err_10 <= w_sys_tmp460;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_alpha_11 <= w_sys_tmp75;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h3b: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_sum_12 <= w_sys_tmp337;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b)) begin
										r_threadTop_sum_12 <= w_sys_tmp340;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b) || (r_sys_threadTop_step==7'h1e) || (r_sys_threadTop_step==7'h21) || (r_sys_threadTop_step==7'h24) || (r_sys_threadTop_step==7'h27)) begin
										r_threadTop_delta_13 <= w_sys_tmp240;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h17) || (r_sys_threadTop_step==7'h19) || (r_sys_threadTop_step==7'h1b) || (r_sys_threadTop_step==7'h1d) || (r_sys_threadTop_step==7'h1f)) begin
										r_threadTop_delta_13 <= w_sys_tmp354;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h7: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_i_14 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h4f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_i_14 <= w_sys_tmp462;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hc: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_15 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_j_15 <= w_sys_tmp87;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h12: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_16 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_16 <= w_sys_tmp180;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_17 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_j_17 <= w_sys_tmp131;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1f: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_18 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_18 <= w_sys_tmp235;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h25: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_19 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_j_19 <= w_sys_tmp194;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h2c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_20 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h2e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_20 <= w_sys_tmp237;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h31: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_21 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_j_21 <= w_sys_tmp258;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h37: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_l_22 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_l_22 <= w_sys_tmp336;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h3d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_23 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_23 <= w_sys_tmp351;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h43: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_j_24 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_j_24 <= w_sys_tmp371;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h4a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_25 <= w_sys_intZero;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_k_25 <= w_sys_tmp459;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'hc: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy0_j_27 <= r_threadTop_j_15;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_copy0_j_27 <= w_sys_tmp86;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h18: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy0_j_28 <= r_threadTop_j_17;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_copy0_j_28 <= w_sys_tmp130;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h25: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy0_j_29 <= r_threadTop_j_19;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_copy0_j_29 <= w_sys_tmp193;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h31: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy0_j_30 <= r_threadTop_j_21;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_copy0_j_30 <= w_sys_tmp256;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h31: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy1_j_31 <= r_threadTop_j_21;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_copy1_j_31 <= w_sys_tmp257;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h43: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy0_j_32 <= r_threadTop_j_24;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_copy0_j_32 <= w_sys_tmp369;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h43: begin

							case(r_sys_threadTop_stage) 
								2'h1: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_threadTop_copy1_j_33 <= r_threadTop_j_24;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h4)) begin
										r_threadTop_copy1_j_33 <= w_sys_tmp370;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1)) begin
										r_sys_tmp0_int <= w_sys_tmp87;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3)) begin
										r_sys_tmp0_int <= w_sys_tmp130;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp0_int <= r_threadTop_k_18;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp0_int <= w_sys_tmp481;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp0_int <= w_sys_tmp488;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp1_int <= r_threadTop_j_15;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp1_int <= w_sys_tmp87;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3)) begin
										r_sys_tmp1_int <= w_sys_tmp471;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp1_int <= w_sys_tmp480;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp1_int <= w_sys_tmp489;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0) || (r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp2_int <= w_sys_tmp87;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp2_int <= r_threadTop_k_16;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3)) begin
										r_sys_tmp2_int <= w_sys_tmp193;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp2_int <= w_sys_tmp481;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp2_int <= w_sys_tmp490;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h10: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3)) begin
										r_sys_tmp3_int <= w_sys_tmp467;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3)) begin
										r_sys_tmp3_int <= w_sys_tmp475;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp3_int <= w_sys_tmp480;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3)) begin
										r_sys_tmp3_int <= w_sys_tmp371;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'ha)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'ha)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_tmp0_float <= w_fld_res_9_dataout_1;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1b)) begin
										r_sys_tmp0_float <= w_sys_tmp354;

									end
									else
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_tmp0_float <= w_fld_input_5_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h9)) begin
										r_sys_tmp1_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h9)) begin
										r_sys_tmp1_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6)) begin
										r_sys_tmp1_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h19)) begin
										r_sys_tmp1_float <= w_sys_tmp354;

									end
									else
									if((r_sys_threadTop_step==7'h5)) begin
										r_sys_tmp1_float <= w_fld_input_5_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_sys_tmp2_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h8)) begin
										r_sys_tmp2_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h5)) begin
										r_sys_tmp2_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1d)) begin
										r_sys_tmp2_float <= w_sys_tmp354;

									end
									else
									if((r_sys_threadTop_step==7'h7) || (r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hb)) begin
										r_sys_tmp2_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_threadTop_step==7'h8) || (r_sys_threadTop_step==7'ha)) begin
										r_sys_tmp2_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h1c: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'hb)) begin
										r_sys_tmp3_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp3_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

						7'h29: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp3_float <= w_fld_output_7_dataout_1;

									end
									else
									if((r_sys_threadTop_step==7'hb)) begin
										r_sys_tmp3_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h4)) begin
										r_sys_tmp3_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1)) begin
										r_sys_tmp4_int <= w_sys_tmp481;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp4_int <= r_threadTop_k_23;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp4_int <= w_sys_tmp489;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1)) begin
										r_sys_tmp5_int <= w_sys_tmp480;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp5_int <= r_threadTop_k_23;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1)) begin
										r_sys_tmp5_int <= w_sys_tmp490;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp6_int <= w_sys_tmp479;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp6_int <= w_sys_tmp490;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp6_int <= r_threadTop_k_25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp7_int <= w_sys_tmp480;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp7_int <= w_sys_tmp489;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp7_int <= w_sys_tmp497;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h0)) begin
										r_sys_tmp8_int <= w_sys_tmp481;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp8_int <= w_sys_tmp490;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((7'h0<=r_sys_threadTop_step && r_sys_threadTop_step<=7'h3)) begin
										r_sys_tmp9_int <= w_sys_tmp258;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1)) begin
										r_sys_tmp9_int <= w_sys_tmp489;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp4_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp4_float <= w_fld_output_7_dataout_1;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3)) begin
										r_sys_tmp4_float <= w_fld_input_5_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp5_float <= w_fld_hidden_6_dataout_1;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h9)) begin
										r_sys_tmp5_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp5_float <= w_fld_w2_4_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp6_float <= w_fld_w2_4_dataout_1;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h4)) begin
										r_sys_tmp6_float <= w_fld_input_5_dataout_1;

									end
								end

							endcase
						end

						7'h4e: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h7)) begin
										r_sys_tmp6_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h6) || (r_sys_threadTop_step==7'hc)) begin
										r_sys_tmp7_float <= w_fld_output_7_dataout_1;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp7_float <= w_fld_input_5_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3) || (r_sys_threadTop_step==7'h5)) begin
										r_sys_tmp8_float <= w_fld_res_9_dataout_1;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h2)) begin
										r_sys_tmp8_float <= w_fld_w1_3_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h3) || (r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hf)) begin
										r_sys_tmp9_float <= w_fld_output_7_dataout_1;

									end
									else
									if((r_sys_threadTop_step==7'h21)) begin
										r_sys_tmp9_float <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_threadTop_phase) 
						7'h35: begin

							case(r_sys_threadTop_stage) 
								2'h0: begin
									if((r_sys_threadTop_step==7'h1e) || (r_sys_threadTop_step==7'h24)) begin
										r_sys_tmp10_float <= w_sys_tmp240;

									end
									else
									if((r_sys_threadTop_step==7'h9) || (r_sys_threadTop_step==7'hc) || (r_sys_threadTop_step==7'hf) || (r_sys_threadTop_step==7'h12) || (r_sys_threadTop_step==7'h15)) begin
										r_sys_tmp10_float <= w_ip_AddFloat_result_0;

									end
									else
									if((r_sys_threadTop_step==7'h4)) begin
										r_sys_tmp10_float <= w_fld_res_9_dataout_1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
