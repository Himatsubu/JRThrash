/*
TimeStamp:	2016/10/27		17:34
*/


module c1(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 9:0] r_sys_run_phase;
	reg         [ 5:0] r_sys_run_stage;
	reg         [ 5:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 5:0] w_sys_run_stage_p1;
	wire        [ 5:0] w_sys_run_step_p1;
	wire signed [14:0] w_fld_u_0_addr_0;
	wire        [31:0] w_fld_u_0_datain_0;
	wire        [31:0] w_fld_u_0_dataout_0;
	wire               w_fld_u_0_r_w_0;
	wire               w_fld_u_0_ce_0;
	reg  signed [14:0] r_fld_u_0_addr_1;
	reg         [31:0] r_fld_u_0_datain_1;
	wire        [31:0] w_fld_u_0_dataout_1;
	reg                r_fld_u_0_r_w_1;
	wire               w_fld_u_0_ce_1;
	reg  signed [31:0] r_run_k_33;
	reg  signed [31:0] r_run_j_34;
	reg  signed [31:0] r_run_n_35;
	reg  signed [31:0] r_run_mx_36;
	reg  signed [31:0] r_run_my_37;
	reg  signed [31:0] r_run_nlast_38;
	reg  signed [31:0] r_run_tmpj_39;
	reg  signed [31:0] r_run_copy0_j_40;
	reg  signed [31:0] r_run_copy0_j_41;
	reg  signed [31:0] r_run_copy0_j_42;
	reg  signed [31:0] r_run_copy0_j_43;
	reg  signed [31:0] r_run_copy0_j_44;
	reg  signed [31:0] r_run_copy0_j_45;
	reg  signed [31:0] r_run_copy0_j_46;
	reg  signed [31:0] r_run_copy0_j_47;
	reg  signed [31:0] r_run_copy0_j_48;
	reg  signed [31:0] r_run_copy0_j_49;
	reg  signed [31:0] r_run_copy0_j_50;
	reg  signed [31:0] r_run_copy0_j_51;
	reg  signed [31:0] r_run_copy0_j_52;
	reg  signed [31:0] r_run_copy0_j_53;
	reg  signed [31:0] r_run_copy0_j_54;
	reg  signed [31:0] r_run_copy0_j_55;
	reg  signed [31:0] r_run_copy0_j_56;
	reg  signed [31:0] r_run_copy0_j_57;
	reg  signed [31:0] r_run_copy0_j_58;
	reg  signed [31:0] r_run_copy0_j_59;
	reg  signed [31:0] r_run_copy0_j_60;
	reg  signed [31:0] r_run_copy0_j_61;
	reg  signed [31:0] r_run_copy0_j_62;
	reg  signed [31:0] r_run_copy0_j_63;
	reg  signed [31:0] r_run_copy0_j_64;
	reg  signed [31:0] r_run_copy0_j_65;
	reg  signed [31:0] r_run_copy0_j_66;
	reg  signed [31:0] r_run_copy0_j_67;
	reg  signed [31:0] r_run_copy0_j_68;
	reg  signed [31:0] r_run_copy0_j_69;
	reg  signed [31:0] r_run_copy0_j_70;
	reg  signed [31:0] r_run_copy0_j_71;
	reg  signed [31:0] r_run_copy0_j_72;
	reg  signed [31:0] r_run_copy1_j_73;
	reg  signed [31:0] r_run_copy2_j_74;
	reg  signed [31:0] r_run_copy3_j_75;
	reg  signed [31:0] r_run_copy4_j_76;
	reg  signed [31:0] r_run_copy5_j_77;
	reg  signed [31:0] r_run_copy6_j_78;
	reg  signed [31:0] r_run_copy7_j_79;
	reg  signed [31:0] r_run_copy8_j_80;
	reg  signed [31:0] r_run_copy9_j_81;
	reg  signed [31:0] r_run_copy10_j_82;
	reg  signed [31:0] r_run_copy0_j_83;
	reg  signed [31:0] r_run_copy1_j_84;
	reg  signed [31:0] r_run_copy2_j_85;
	reg  signed [31:0] r_run_copy3_j_86;
	reg  signed [31:0] r_run_copy4_j_87;
	reg  signed [31:0] r_run_copy5_j_88;
	reg  signed [31:0] r_run_copy6_j_89;
	reg  signed [31:0] r_run_copy7_j_90;
	reg  signed [31:0] r_run_copy8_j_91;
	reg  signed [31:0] r_run_copy9_j_92;
	reg  signed [31:0] r_run_copy10_j_93;
	reg  signed [31:0] r_run_copy0_j_94;
	reg  signed [31:0] r_run_copy1_j_95;
	reg  signed [31:0] r_run_copy2_j_96;
	reg  signed [31:0] r_run_copy3_j_97;
	reg  signed [31:0] r_run_copy4_j_98;
	reg  signed [31:0] r_run_copy5_j_99;
	reg  signed [31:0] r_run_copy6_j_100;
	reg  signed [31:0] r_run_copy7_j_101;
	reg  signed [31:0] r_run_copy8_j_102;
	reg  signed [31:0] r_run_copy9_j_103;
	reg  signed [31:0] r_run_copy10_j_104;
	reg  signed [31:0] r_run_copy0_j_105;
	reg  signed [31:0] r_run_copy1_j_106;
	reg  signed [31:0] r_run_copy2_j_107;
	reg  signed [31:0] r_run_copy3_j_108;
	reg  signed [31:0] r_run_copy4_j_109;
	reg  signed [31:0] r_run_copy5_j_110;
	reg  signed [31:0] r_run_copy6_j_111;
	reg  signed [31:0] r_run_copy7_j_112;
	reg  signed [31:0] r_run_copy8_j_113;
	reg  signed [31:0] r_run_copy9_j_114;
	reg  signed [31:0] r_run_copy10_j_115;
	reg  signed [31:0] r_run_copy0_j_116;
	reg  signed [31:0] r_run_copy1_j_117;
	reg  signed [31:0] r_run_copy2_j_118;
	reg  signed [31:0] r_run_copy3_j_119;
	reg  signed [31:0] r_run_copy4_j_120;
	reg  signed [31:0] r_run_copy5_j_121;
	reg  signed [31:0] r_run_copy6_j_122;
	reg  signed [31:0] r_run_copy7_j_123;
	reg  signed [31:0] r_run_copy8_j_124;
	reg  signed [31:0] r_run_copy9_j_125;
	reg  signed [31:0] r_run_copy10_j_126;
	reg  signed [31:0] r_run_copy0_j_127;
	reg  signed [31:0] r_run_copy1_j_128;
	reg  signed [31:0] r_run_copy2_j_129;
	reg  signed [31:0] r_run_copy3_j_130;
	reg  signed [31:0] r_run_copy4_j_131;
	reg  signed [31:0] r_run_copy5_j_132;
	reg  signed [31:0] r_run_copy6_j_133;
	reg  signed [31:0] r_run_copy7_j_134;
	reg  signed [31:0] r_run_copy8_j_135;
	reg  signed [31:0] r_run_copy9_j_136;
	reg  signed [31:0] r_run_copy10_j_137;
	reg  signed [31:0] r_run_copy0_j_138;
	reg  signed [31:0] r_run_copy1_j_139;
	reg  signed [31:0] r_run_copy2_j_140;
	reg  signed [31:0] r_run_copy3_j_141;
	reg  signed [31:0] r_run_copy4_j_142;
	reg  signed [31:0] r_run_copy5_j_143;
	reg  signed [31:0] r_run_copy6_j_144;
	reg  signed [31:0] r_run_copy7_j_145;
	reg  signed [31:0] r_run_copy8_j_146;
	reg  signed [31:0] r_run_copy9_j_147;
	reg  signed [31:0] r_run_copy10_j_148;
	reg  signed [31:0] r_run_copy0_j_149;
	reg  signed [31:0] r_run_copy1_j_150;
	reg  signed [31:0] r_run_copy2_j_151;
	reg  signed [31:0] r_run_copy3_j_152;
	reg  signed [31:0] r_run_copy4_j_153;
	reg  signed [31:0] r_run_copy5_j_154;
	reg  signed [31:0] r_run_copy6_j_155;
	reg  signed [31:0] r_run_copy7_j_156;
	reg  signed [31:0] r_run_copy8_j_157;
	reg  signed [31:0] r_run_copy9_j_158;
	reg  signed [31:0] r_run_copy10_j_159;
	reg  signed [31:0] r_run_copy0_j_160;
	reg  signed [31:0] r_run_copy0_j_161;
	reg  signed [31:0] r_run_copy1_j_162;
	reg  signed [31:0] r_run_copy0_j_163;
	reg  signed [31:0] r_run_copy1_j_164;
	reg  signed [31:0] r_run_copy0_j_165;
	reg  signed [31:0] r_run_copy1_j_166;
	reg  signed [31:0] r_run_copy0_j_167;
	reg  signed [31:0] r_run_copy1_j_168;
	reg  signed [31:0] r_run_copy0_j_169;
	reg  signed [31:0] r_run_copy1_j_170;
	reg  signed [31:0] r_run_copy0_j_171;
	reg  signed [31:0] r_run_copy1_j_172;
	reg  signed [31:0] r_run_copy0_j_173;
	reg  signed [31:0] r_run_copy1_j_174;
	reg  signed [31:0] r_run_copy0_j_175;
	reg  signed [31:0] r_run_copy0_j_176;
	reg  signed [31:0] r_run_copy1_j_177;
	reg  signed [31:0] r_run_copy0_j_178;
	reg  signed [31:0] r_run_copy1_j_179;
	reg  signed [31:0] r_run_copy0_j_180;
	reg  signed [31:0] r_run_copy1_j_181;
	reg  signed [31:0] r_run_copy0_j_182;
	reg  signed [31:0] r_run_copy1_j_183;
	reg  signed [31:0] r_run_copy0_j_184;
	reg  signed [31:0] r_run_copy1_j_185;
	reg  signed [31:0] r_run_copy0_j_186;
	reg  signed [31:0] r_run_copy1_j_187;
	reg  signed [31:0] r_run_copy0_j_188;
	reg  signed [31:0] r_run_copy1_j_189;
	reg  signed [31:0] r_run_copy0_j_190;
	reg  signed [31:0] r_run_copy0_j_191;
	reg  signed [31:0] r_run_copy1_j_192;
	reg  signed [31:0] r_run_copy0_j_193;
	reg  signed [31:0] r_run_copy1_j_194;
	reg  signed [31:0] r_run_copy0_j_195;
	reg  signed [31:0] r_run_copy1_j_196;
	reg  signed [31:0] r_run_copy0_j_197;
	reg  signed [31:0] r_run_copy1_j_198;
	reg  signed [31:0] r_run_copy0_j_199;
	reg  signed [31:0] r_run_copy1_j_200;
	reg  signed [31:0] r_run_copy0_j_201;
	reg  signed [31:0] r_run_copy1_j_202;
	reg  signed [31:0] r_run_copy0_j_203;
	reg  signed [31:0] r_run_copy1_j_204;
	reg  signed [31:0] r_run_copy0_j_205;
	reg  signed [31:0] r_run_copy0_j_206;
	reg  signed [31:0] r_run_copy1_j_207;
	reg  signed [31:0] r_run_copy0_j_208;
	reg  signed [31:0] r_run_copy1_j_209;
	reg  signed [31:0] r_run_copy0_j_210;
	reg  signed [31:0] r_run_copy1_j_211;
	reg  signed [31:0] r_run_copy0_j_212;
	reg  signed [31:0] r_run_copy1_j_213;
	reg  signed [31:0] r_run_copy0_j_214;
	reg  signed [31:0] r_run_copy1_j_215;
	reg  signed [31:0] r_run_copy0_j_216;
	reg  signed [31:0] r_run_copy1_j_217;
	reg  signed [31:0] r_run_copy0_j_218;
	reg  signed [31:0] r_run_copy1_j_219;
	reg                r_sub19_run_req;
	wire               w_sub19_run_busy;
	wire signed [11:0] w_sub19_u_addr;
	reg  signed [11:0] r_sub19_u_addr;
	wire        [31:0] w_sub19_u_datain;
	reg         [31:0] r_sub19_u_datain;
	wire        [31:0] w_sub19_u_dataout;
	wire               w_sub19_u_r_w;
	reg                r_sub19_u_r_w;
	wire signed [11:0] w_sub19_result_addr;
	reg  signed [11:0] r_sub19_result_addr;
	wire        [31:0] w_sub19_result_datain;
	reg         [31:0] r_sub19_result_datain;
	wire        [31:0] w_sub19_result_dataout;
	wire               w_sub19_result_r_w;
	reg                r_sub19_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [11:0] w_sub12_u_addr;
	reg  signed [11:0] r_sub12_u_addr;
	wire        [31:0] w_sub12_u_datain;
	reg         [31:0] r_sub12_u_datain;
	wire        [31:0] w_sub12_u_dataout;
	wire               w_sub12_u_r_w;
	reg                r_sub12_u_r_w;
	wire signed [11:0] w_sub12_result_addr;
	reg  signed [11:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [11:0] w_sub11_u_addr;
	reg  signed [11:0] r_sub11_u_addr;
	wire        [31:0] w_sub11_u_datain;
	reg         [31:0] r_sub11_u_datain;
	wire        [31:0] w_sub11_u_dataout;
	wire               w_sub11_u_r_w;
	reg                r_sub11_u_r_w;
	wire signed [11:0] w_sub11_result_addr;
	reg  signed [11:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [11:0] w_sub14_u_addr;
	reg  signed [11:0] r_sub14_u_addr;
	wire        [31:0] w_sub14_u_datain;
	reg         [31:0] r_sub14_u_datain;
	wire        [31:0] w_sub14_u_dataout;
	wire               w_sub14_u_r_w;
	reg                r_sub14_u_r_w;
	wire signed [11:0] w_sub14_result_addr;
	reg  signed [11:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [11:0] w_sub13_u_addr;
	reg  signed [11:0] r_sub13_u_addr;
	wire        [31:0] w_sub13_u_datain;
	reg         [31:0] r_sub13_u_datain;
	wire        [31:0] w_sub13_u_dataout;
	wire               w_sub13_u_r_w;
	reg                r_sub13_u_r_w;
	wire signed [11:0] w_sub13_result_addr;
	reg  signed [11:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub16_run_req;
	wire               w_sub16_run_busy;
	wire signed [11:0] w_sub16_u_addr;
	reg  signed [11:0] r_sub16_u_addr;
	wire        [31:0] w_sub16_u_datain;
	reg         [31:0] r_sub16_u_datain;
	wire        [31:0] w_sub16_u_dataout;
	wire               w_sub16_u_r_w;
	reg                r_sub16_u_r_w;
	wire signed [11:0] w_sub16_result_addr;
	reg  signed [11:0] r_sub16_result_addr;
	wire        [31:0] w_sub16_result_datain;
	reg         [31:0] r_sub16_result_datain;
	wire        [31:0] w_sub16_result_dataout;
	wire               w_sub16_result_r_w;
	reg                r_sub16_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [11:0] w_sub15_u_addr;
	reg  signed [11:0] r_sub15_u_addr;
	wire        [31:0] w_sub15_u_datain;
	reg         [31:0] r_sub15_u_datain;
	wire        [31:0] w_sub15_u_dataout;
	wire               w_sub15_u_r_w;
	reg                r_sub15_u_r_w;
	wire signed [11:0] w_sub15_result_addr;
	reg  signed [11:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub18_run_req;
	wire               w_sub18_run_busy;
	wire signed [11:0] w_sub18_u_addr;
	reg  signed [11:0] r_sub18_u_addr;
	wire        [31:0] w_sub18_u_datain;
	reg         [31:0] r_sub18_u_datain;
	wire        [31:0] w_sub18_u_dataout;
	wire               w_sub18_u_r_w;
	reg                r_sub18_u_r_w;
	wire signed [11:0] w_sub18_result_addr;
	reg  signed [11:0] r_sub18_result_addr;
	wire        [31:0] w_sub18_result_datain;
	reg         [31:0] r_sub18_result_datain;
	wire        [31:0] w_sub18_result_dataout;
	wire               w_sub18_result_r_w;
	reg                r_sub18_result_r_w;
	reg                r_sub17_run_req;
	wire               w_sub17_run_busy;
	wire signed [11:0] w_sub17_u_addr;
	reg  signed [11:0] r_sub17_u_addr;
	wire        [31:0] w_sub17_u_datain;
	reg         [31:0] r_sub17_u_datain;
	wire        [31:0] w_sub17_u_dataout;
	wire               w_sub17_u_r_w;
	reg                r_sub17_u_r_w;
	wire signed [11:0] w_sub17_result_addr;
	reg  signed [11:0] r_sub17_result_addr;
	wire        [31:0] w_sub17_result_datain;
	reg         [31:0] r_sub17_result_datain;
	wire        [31:0] w_sub17_result_dataout;
	wire               w_sub17_result_r_w;
	reg                r_sub17_result_r_w;
	reg                r_sub20_run_req;
	wire               w_sub20_run_busy;
	wire signed [11:0] w_sub20_u_addr;
	reg  signed [11:0] r_sub20_u_addr;
	wire        [31:0] w_sub20_u_datain;
	reg         [31:0] r_sub20_u_datain;
	wire        [31:0] w_sub20_u_dataout;
	wire               w_sub20_u_r_w;
	reg                r_sub20_u_r_w;
	wire signed [11:0] w_sub20_result_addr;
	reg  signed [11:0] r_sub20_result_addr;
	wire        [31:0] w_sub20_result_datain;
	reg         [31:0] r_sub20_result_datain;
	wire        [31:0] w_sub20_result_dataout;
	wire               w_sub20_result_r_w;
	reg                r_sub20_result_r_w;
	reg                r_sub21_run_req;
	wire               w_sub21_run_busy;
	wire signed [11:0] w_sub21_u_addr;
	reg  signed [11:0] r_sub21_u_addr;
	wire        [31:0] w_sub21_u_datain;
	reg         [31:0] r_sub21_u_datain;
	wire        [31:0] w_sub21_u_dataout;
	wire               w_sub21_u_r_w;
	reg                r_sub21_u_r_w;
	wire signed [11:0] w_sub21_result_addr;
	reg  signed [11:0] r_sub21_result_addr;
	wire        [31:0] w_sub21_result_datain;
	reg         [31:0] r_sub21_result_datain;
	wire        [31:0] w_sub21_result_dataout;
	wire               w_sub21_result_r_w;
	reg                r_sub21_result_r_w;
	reg                r_sub28_run_req;
	wire               w_sub28_run_busy;
	wire signed [11:0] w_sub28_u_addr;
	reg  signed [11:0] r_sub28_u_addr;
	wire        [31:0] w_sub28_u_datain;
	reg         [31:0] r_sub28_u_datain;
	wire        [31:0] w_sub28_u_dataout;
	wire               w_sub28_u_r_w;
	reg                r_sub28_u_r_w;
	wire signed [11:0] w_sub28_result_addr;
	reg  signed [11:0] r_sub28_result_addr;
	wire        [31:0] w_sub28_result_datain;
	reg         [31:0] r_sub28_result_datain;
	wire        [31:0] w_sub28_result_dataout;
	wire               w_sub28_result_r_w;
	reg                r_sub28_result_r_w;
	reg                r_sub29_run_req;
	wire               w_sub29_run_busy;
	wire signed [11:0] w_sub29_u_addr;
	reg  signed [11:0] r_sub29_u_addr;
	wire        [31:0] w_sub29_u_datain;
	reg         [31:0] r_sub29_u_datain;
	wire        [31:0] w_sub29_u_dataout;
	wire               w_sub29_u_r_w;
	reg                r_sub29_u_r_w;
	wire signed [11:0] w_sub29_result_addr;
	reg  signed [11:0] r_sub29_result_addr;
	wire        [31:0] w_sub29_result_datain;
	reg         [31:0] r_sub29_result_datain;
	wire        [31:0] w_sub29_result_dataout;
	wire               w_sub29_result_r_w;
	reg                r_sub29_result_r_w;
	reg                r_sub26_run_req;
	wire               w_sub26_run_busy;
	wire signed [11:0] w_sub26_u_addr;
	reg  signed [11:0] r_sub26_u_addr;
	wire        [31:0] w_sub26_u_datain;
	reg         [31:0] r_sub26_u_datain;
	wire        [31:0] w_sub26_u_dataout;
	wire               w_sub26_u_r_w;
	reg                r_sub26_u_r_w;
	wire signed [11:0] w_sub26_result_addr;
	reg  signed [11:0] r_sub26_result_addr;
	wire        [31:0] w_sub26_result_datain;
	reg         [31:0] r_sub26_result_datain;
	wire        [31:0] w_sub26_result_dataout;
	wire               w_sub26_result_r_w;
	reg                r_sub26_result_r_w;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [11:0] w_sub09_u_addr;
	reg  signed [11:0] r_sub09_u_addr;
	wire        [31:0] w_sub09_u_datain;
	reg         [31:0] r_sub09_u_datain;
	wire        [31:0] w_sub09_u_dataout;
	wire               w_sub09_u_r_w;
	reg                r_sub09_u_r_w;
	wire signed [11:0] w_sub09_result_addr;
	reg  signed [11:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub27_run_req;
	wire               w_sub27_run_busy;
	wire signed [11:0] w_sub27_u_addr;
	reg  signed [11:0] r_sub27_u_addr;
	wire        [31:0] w_sub27_u_datain;
	reg         [31:0] r_sub27_u_datain;
	wire        [31:0] w_sub27_u_dataout;
	wire               w_sub27_u_r_w;
	reg                r_sub27_u_r_w;
	wire signed [11:0] w_sub27_result_addr;
	reg  signed [11:0] r_sub27_result_addr;
	wire        [31:0] w_sub27_result_datain;
	reg         [31:0] r_sub27_result_datain;
	wire        [31:0] w_sub27_result_dataout;
	wire               w_sub27_result_r_w;
	reg                r_sub27_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [11:0] w_sub08_u_addr;
	reg  signed [11:0] r_sub08_u_addr;
	wire        [31:0] w_sub08_u_datain;
	reg         [31:0] r_sub08_u_datain;
	wire        [31:0] w_sub08_u_dataout;
	wire               w_sub08_u_r_w;
	reg                r_sub08_u_r_w;
	wire signed [11:0] w_sub08_result_addr;
	reg  signed [11:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub24_run_req;
	wire               w_sub24_run_busy;
	wire signed [11:0] w_sub24_u_addr;
	reg  signed [11:0] r_sub24_u_addr;
	wire        [31:0] w_sub24_u_datain;
	reg         [31:0] r_sub24_u_datain;
	wire        [31:0] w_sub24_u_dataout;
	wire               w_sub24_u_r_w;
	reg                r_sub24_u_r_w;
	wire signed [11:0] w_sub24_result_addr;
	reg  signed [11:0] r_sub24_result_addr;
	wire        [31:0] w_sub24_result_datain;
	reg         [31:0] r_sub24_result_datain;
	wire        [31:0] w_sub24_result_dataout;
	wire               w_sub24_result_r_w;
	reg                r_sub24_result_r_w;
	reg                r_sub25_run_req;
	wire               w_sub25_run_busy;
	wire signed [11:0] w_sub25_u_addr;
	reg  signed [11:0] r_sub25_u_addr;
	wire        [31:0] w_sub25_u_datain;
	reg         [31:0] r_sub25_u_datain;
	wire        [31:0] w_sub25_u_dataout;
	wire               w_sub25_u_r_w;
	reg                r_sub25_u_r_w;
	wire signed [11:0] w_sub25_result_addr;
	reg  signed [11:0] r_sub25_result_addr;
	wire        [31:0] w_sub25_result_datain;
	reg         [31:0] r_sub25_result_datain;
	wire        [31:0] w_sub25_result_dataout;
	wire               w_sub25_result_r_w;
	reg                r_sub25_result_r_w;
	reg                r_sub22_run_req;
	wire               w_sub22_run_busy;
	wire signed [11:0] w_sub22_u_addr;
	reg  signed [11:0] r_sub22_u_addr;
	wire        [31:0] w_sub22_u_datain;
	reg         [31:0] r_sub22_u_datain;
	wire        [31:0] w_sub22_u_dataout;
	wire               w_sub22_u_r_w;
	reg                r_sub22_u_r_w;
	wire signed [11:0] w_sub22_result_addr;
	reg  signed [11:0] r_sub22_result_addr;
	wire        [31:0] w_sub22_result_datain;
	reg         [31:0] r_sub22_result_datain;
	wire        [31:0] w_sub22_result_dataout;
	wire               w_sub22_result_r_w;
	reg                r_sub22_result_r_w;
	reg                r_sub23_run_req;
	wire               w_sub23_run_busy;
	wire signed [11:0] w_sub23_u_addr;
	reg  signed [11:0] r_sub23_u_addr;
	wire        [31:0] w_sub23_u_datain;
	reg         [31:0] r_sub23_u_datain;
	wire        [31:0] w_sub23_u_dataout;
	wire               w_sub23_u_r_w;
	reg                r_sub23_u_r_w;
	wire signed [11:0] w_sub23_result_addr;
	reg  signed [11:0] r_sub23_result_addr;
	wire        [31:0] w_sub23_result_datain;
	reg         [31:0] r_sub23_result_datain;
	wire        [31:0] w_sub23_result_dataout;
	wire               w_sub23_result_r_w;
	reg                r_sub23_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [11:0] w_sub03_u_addr;
	reg  signed [11:0] r_sub03_u_addr;
	wire        [31:0] w_sub03_u_datain;
	reg         [31:0] r_sub03_u_datain;
	wire        [31:0] w_sub03_u_dataout;
	wire               w_sub03_u_r_w;
	reg                r_sub03_u_r_w;
	wire signed [11:0] w_sub03_result_addr;
	reg  signed [11:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [11:0] w_sub02_u_addr;
	reg  signed [11:0] r_sub02_u_addr;
	wire        [31:0] w_sub02_u_datain;
	reg         [31:0] r_sub02_u_datain;
	wire        [31:0] w_sub02_u_dataout;
	wire               w_sub02_u_r_w;
	reg                r_sub02_u_r_w;
	wire signed [11:0] w_sub02_result_addr;
	reg  signed [11:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [11:0] w_sub01_u_addr;
	reg  signed [11:0] r_sub01_u_addr;
	wire        [31:0] w_sub01_u_datain;
	reg         [31:0] r_sub01_u_datain;
	wire        [31:0] w_sub01_u_dataout;
	wire               w_sub01_u_r_w;
	reg                r_sub01_u_r_w;
	wire signed [11:0] w_sub01_result_addr;
	reg  signed [11:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [11:0] w_sub00_u_addr;
	reg  signed [11:0] r_sub00_u_addr;
	wire        [31:0] w_sub00_u_datain;
	reg         [31:0] r_sub00_u_datain;
	wire        [31:0] w_sub00_u_dataout;
	wire               w_sub00_u_r_w;
	reg                r_sub00_u_r_w;
	wire signed [11:0] w_sub00_result_addr;
	reg  signed [11:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [11:0] w_sub07_u_addr;
	reg  signed [11:0] r_sub07_u_addr;
	wire        [31:0] w_sub07_u_datain;
	reg         [31:0] r_sub07_u_datain;
	wire        [31:0] w_sub07_u_dataout;
	wire               w_sub07_u_r_w;
	reg                r_sub07_u_r_w;
	wire signed [11:0] w_sub07_result_addr;
	reg  signed [11:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [11:0] w_sub06_u_addr;
	reg  signed [11:0] r_sub06_u_addr;
	wire        [31:0] w_sub06_u_datain;
	reg         [31:0] r_sub06_u_datain;
	wire        [31:0] w_sub06_u_dataout;
	wire               w_sub06_u_r_w;
	reg                r_sub06_u_r_w;
	wire signed [11:0] w_sub06_result_addr;
	reg  signed [11:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [11:0] w_sub05_u_addr;
	reg  signed [11:0] r_sub05_u_addr;
	wire        [31:0] w_sub05_u_datain;
	reg         [31:0] r_sub05_u_datain;
	wire        [31:0] w_sub05_u_dataout;
	wire               w_sub05_u_r_w;
	reg                r_sub05_u_r_w;
	wire signed [11:0] w_sub05_result_addr;
	reg  signed [11:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [11:0] w_sub04_u_addr;
	reg  signed [11:0] r_sub04_u_addr;
	wire        [31:0] w_sub04_u_datain;
	reg         [31:0] r_sub04_u_datain;
	wire        [31:0] w_sub04_u_dataout;
	wire               w_sub04_u_r_w;
	reg                r_sub04_u_r_w;
	wire signed [11:0] w_sub04_result_addr;
	reg  signed [11:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [11:0] w_sub10_u_addr;
	reg  signed [11:0] r_sub10_u_addr;
	wire        [31:0] w_sub10_u_datain;
	reg         [31:0] r_sub10_u_datain;
	wire        [31:0] w_sub10_u_dataout;
	wire               w_sub10_u_r_w;
	reg                r_sub10_u_r_w;
	wire signed [11:0] w_sub10_result_addr;
	reg  signed [11:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg                r_sub31_run_req;
	wire               w_sub31_run_busy;
	wire signed [11:0] w_sub31_u_addr;
	reg  signed [11:0] r_sub31_u_addr;
	wire        [31:0] w_sub31_u_datain;
	reg         [31:0] r_sub31_u_datain;
	wire        [31:0] w_sub31_u_dataout;
	wire               w_sub31_u_r_w;
	reg                r_sub31_u_r_w;
	wire signed [11:0] w_sub31_result_addr;
	reg  signed [11:0] r_sub31_result_addr;
	wire        [31:0] w_sub31_result_datain;
	reg         [31:0] r_sub31_result_datain;
	wire        [31:0] w_sub31_result_dataout;
	wire               w_sub31_result_r_w;
	reg                r_sub31_result_r_w;
	reg                r_sub30_run_req;
	wire               w_sub30_run_busy;
	wire signed [11:0] w_sub30_u_addr;
	reg  signed [11:0] r_sub30_u_addr;
	wire        [31:0] w_sub30_u_datain;
	reg         [31:0] r_sub30_u_datain;
	wire        [31:0] w_sub30_u_dataout;
	wire               w_sub30_u_r_w;
	reg                r_sub30_u_r_w;
	wire signed [11:0] w_sub30_result_addr;
	reg  signed [11:0] r_sub30_result_addr;
	wire        [31:0] w_sub30_result_datain;
	reg         [31:0] r_sub30_result_datain;
	wire        [31:0] w_sub30_result_dataout;
	wire               w_sub30_result_r_w;
	reg                r_sub30_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	wire signed [31:0] w_sys_tmp1;
	wire               w_sys_tmp3;
	wire               w_sys_tmp4;
	wire signed [31:0] w_sys_tmp5;
	wire               w_sys_tmp6;
	wire               w_sys_tmp7;
	wire signed [31:0] w_sys_tmp10;
	wire signed [31:0] w_sys_tmp11;
	wire signed [31:0] w_sys_tmp12;
	wire        [31:0] w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp51;
	wire               w_sys_tmp52;
	wire signed [31:0] w_sys_tmp53;
	wire signed [31:0] w_sys_tmp54;
	wire               w_sys_tmp55;
	wire               w_sys_tmp56;
	wire signed [31:0] w_sys_tmp57;
	wire signed [31:0] w_sys_tmp60;
	wire signed [31:0] w_sys_tmp61;
	wire signed [31:0] w_sys_tmp62;
	wire        [31:0] w_sys_tmp63;
	wire signed [31:0] w_sys_tmp64;
	wire signed [31:0] w_sys_tmp65;
	wire signed [31:0] w_sys_tmp67;
	wire signed [31:0] w_sys_tmp68;
	wire signed [31:0] w_sys_tmp129;
	wire               w_sys_tmp130;
	wire               w_sys_tmp131;
	wire signed [31:0] w_sys_tmp132;
	wire signed [31:0] w_sys_tmp134;
	wire signed [31:0] w_sys_tmp135;
	wire signed [31:0] w_sys_tmp137;
	wire signed [31:0] w_sys_tmp138;
	wire signed [31:0] w_sys_tmp139;
	wire        [31:0] w_sys_tmp140;
	wire signed [31:0] w_sys_tmp141;
	wire signed [31:0] w_sys_tmp142;
	wire signed [31:0] w_sys_tmp144;
	wire signed [31:0] w_sys_tmp145;
	wire signed [31:0] w_sys_tmp218;
	wire               w_sys_tmp219;
	wire               w_sys_tmp220;
	wire signed [31:0] w_sys_tmp221;
	wire signed [31:0] w_sys_tmp223;
	wire signed [31:0] w_sys_tmp224;
	wire signed [31:0] w_sys_tmp226;
	wire signed [31:0] w_sys_tmp227;
	wire signed [31:0] w_sys_tmp228;
	wire        [31:0] w_sys_tmp229;
	wire signed [31:0] w_sys_tmp230;
	wire signed [31:0] w_sys_tmp231;
	wire signed [31:0] w_sys_tmp233;
	wire signed [31:0] w_sys_tmp234;
	wire signed [31:0] w_sys_tmp307;
	wire               w_sys_tmp308;
	wire               w_sys_tmp309;
	wire signed [31:0] w_sys_tmp310;
	wire signed [31:0] w_sys_tmp312;
	wire signed [31:0] w_sys_tmp313;
	wire signed [31:0] w_sys_tmp315;
	wire signed [31:0] w_sys_tmp316;
	wire signed [31:0] w_sys_tmp317;
	wire        [31:0] w_sys_tmp318;
	wire signed [31:0] w_sys_tmp319;
	wire signed [31:0] w_sys_tmp320;
	wire signed [31:0] w_sys_tmp322;
	wire signed [31:0] w_sys_tmp323;
	wire signed [31:0] w_sys_tmp396;
	wire               w_sys_tmp397;
	wire               w_sys_tmp398;
	wire signed [31:0] w_sys_tmp399;
	wire signed [31:0] w_sys_tmp401;
	wire signed [31:0] w_sys_tmp402;
	wire signed [31:0] w_sys_tmp404;
	wire signed [31:0] w_sys_tmp405;
	wire signed [31:0] w_sys_tmp406;
	wire        [31:0] w_sys_tmp407;
	wire signed [31:0] w_sys_tmp408;
	wire signed [31:0] w_sys_tmp409;
	wire signed [31:0] w_sys_tmp411;
	wire signed [31:0] w_sys_tmp412;
	wire signed [31:0] w_sys_tmp485;
	wire               w_sys_tmp486;
	wire               w_sys_tmp487;
	wire signed [31:0] w_sys_tmp488;
	wire signed [31:0] w_sys_tmp490;
	wire signed [31:0] w_sys_tmp491;
	wire signed [31:0] w_sys_tmp493;
	wire signed [31:0] w_sys_tmp494;
	wire signed [31:0] w_sys_tmp495;
	wire        [31:0] w_sys_tmp496;
	wire signed [31:0] w_sys_tmp497;
	wire signed [31:0] w_sys_tmp498;
	wire signed [31:0] w_sys_tmp500;
	wire signed [31:0] w_sys_tmp501;
	wire signed [31:0] w_sys_tmp574;
	wire               w_sys_tmp575;
	wire               w_sys_tmp576;
	wire signed [31:0] w_sys_tmp577;
	wire signed [31:0] w_sys_tmp579;
	wire signed [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp582;
	wire signed [31:0] w_sys_tmp583;
	wire signed [31:0] w_sys_tmp584;
	wire        [31:0] w_sys_tmp585;
	wire signed [31:0] w_sys_tmp586;
	wire signed [31:0] w_sys_tmp587;
	wire signed [31:0] w_sys_tmp589;
	wire signed [31:0] w_sys_tmp590;
	wire signed [31:0] w_sys_tmp663;
	wire               w_sys_tmp664;
	wire               w_sys_tmp665;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp668;
	wire signed [31:0] w_sys_tmp669;
	wire signed [31:0] w_sys_tmp671;
	wire signed [31:0] w_sys_tmp672;
	wire signed [31:0] w_sys_tmp673;
	wire        [31:0] w_sys_tmp674;
	wire signed [31:0] w_sys_tmp675;
	wire signed [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp678;
	wire signed [31:0] w_sys_tmp679;
	wire signed [31:0] w_sys_tmp752;
	wire               w_sys_tmp753;
	wire               w_sys_tmp754;
	wire signed [31:0] w_sys_tmp755;
	wire signed [31:0] w_sys_tmp756;
	wire               w_sys_tmp757;
	wire               w_sys_tmp758;
	wire signed [31:0] w_sys_tmp759;
	wire signed [31:0] w_sys_tmp762;
	wire signed [31:0] w_sys_tmp763;
	wire signed [31:0] w_sys_tmp764;
	wire        [31:0] w_sys_tmp765;
	wire signed [31:0] w_sys_tmp766;
	wire signed [31:0] w_sys_tmp767;
	wire signed [31:0] w_sys_tmp769;
	wire signed [31:0] w_sys_tmp770;
	wire signed [31:0] w_sys_tmp831;
	wire               w_sys_tmp832;
	wire               w_sys_tmp833;
	wire signed [31:0] w_sys_tmp834;
	wire signed [31:0] w_sys_tmp836;
	wire signed [31:0] w_sys_tmp837;
	wire signed [31:0] w_sys_tmp839;
	wire signed [31:0] w_sys_tmp840;
	wire signed [31:0] w_sys_tmp841;
	wire        [31:0] w_sys_tmp842;
	wire signed [31:0] w_sys_tmp843;
	wire signed [31:0] w_sys_tmp844;
	wire signed [31:0] w_sys_tmp846;
	wire signed [31:0] w_sys_tmp847;
	wire signed [31:0] w_sys_tmp920;
	wire               w_sys_tmp921;
	wire               w_sys_tmp922;
	wire signed [31:0] w_sys_tmp923;
	wire signed [31:0] w_sys_tmp925;
	wire signed [31:0] w_sys_tmp926;
	wire signed [31:0] w_sys_tmp928;
	wire signed [31:0] w_sys_tmp929;
	wire signed [31:0] w_sys_tmp930;
	wire        [31:0] w_sys_tmp931;
	wire signed [31:0] w_sys_tmp932;
	wire signed [31:0] w_sys_tmp933;
	wire signed [31:0] w_sys_tmp935;
	wire signed [31:0] w_sys_tmp936;
	wire signed [31:0] w_sys_tmp1009;
	wire               w_sys_tmp1010;
	wire               w_sys_tmp1011;
	wire signed [31:0] w_sys_tmp1012;
	wire signed [31:0] w_sys_tmp1014;
	wire signed [31:0] w_sys_tmp1015;
	wire signed [31:0] w_sys_tmp1017;
	wire signed [31:0] w_sys_tmp1018;
	wire signed [31:0] w_sys_tmp1019;
	wire        [31:0] w_sys_tmp1020;
	wire signed [31:0] w_sys_tmp1021;
	wire signed [31:0] w_sys_tmp1022;
	wire signed [31:0] w_sys_tmp1024;
	wire signed [31:0] w_sys_tmp1025;
	wire signed [31:0] w_sys_tmp1098;
	wire               w_sys_tmp1099;
	wire               w_sys_tmp1100;
	wire signed [31:0] w_sys_tmp1101;
	wire signed [31:0] w_sys_tmp1103;
	wire signed [31:0] w_sys_tmp1104;
	wire signed [31:0] w_sys_tmp1106;
	wire signed [31:0] w_sys_tmp1107;
	wire signed [31:0] w_sys_tmp1108;
	wire        [31:0] w_sys_tmp1109;
	wire signed [31:0] w_sys_tmp1110;
	wire signed [31:0] w_sys_tmp1111;
	wire signed [31:0] w_sys_tmp1113;
	wire signed [31:0] w_sys_tmp1114;
	wire signed [31:0] w_sys_tmp1187;
	wire               w_sys_tmp1188;
	wire               w_sys_tmp1189;
	wire signed [31:0] w_sys_tmp1190;
	wire signed [31:0] w_sys_tmp1192;
	wire signed [31:0] w_sys_tmp1193;
	wire signed [31:0] w_sys_tmp1195;
	wire signed [31:0] w_sys_tmp1196;
	wire signed [31:0] w_sys_tmp1197;
	wire        [31:0] w_sys_tmp1198;
	wire signed [31:0] w_sys_tmp1199;
	wire signed [31:0] w_sys_tmp1200;
	wire signed [31:0] w_sys_tmp1202;
	wire signed [31:0] w_sys_tmp1203;
	wire signed [31:0] w_sys_tmp1276;
	wire               w_sys_tmp1277;
	wire               w_sys_tmp1278;
	wire signed [31:0] w_sys_tmp1279;
	wire signed [31:0] w_sys_tmp1281;
	wire signed [31:0] w_sys_tmp1282;
	wire signed [31:0] w_sys_tmp1284;
	wire signed [31:0] w_sys_tmp1285;
	wire signed [31:0] w_sys_tmp1286;
	wire        [31:0] w_sys_tmp1287;
	wire signed [31:0] w_sys_tmp1288;
	wire signed [31:0] w_sys_tmp1289;
	wire signed [31:0] w_sys_tmp1291;
	wire signed [31:0] w_sys_tmp1292;
	wire signed [31:0] w_sys_tmp1365;
	wire               w_sys_tmp1366;
	wire               w_sys_tmp1367;
	wire signed [31:0] w_sys_tmp1368;
	wire signed [31:0] w_sys_tmp1370;
	wire signed [31:0] w_sys_tmp1371;
	wire signed [31:0] w_sys_tmp1373;
	wire signed [31:0] w_sys_tmp1374;
	wire signed [31:0] w_sys_tmp1375;
	wire        [31:0] w_sys_tmp1376;
	wire signed [31:0] w_sys_tmp1377;
	wire signed [31:0] w_sys_tmp1378;
	wire signed [31:0] w_sys_tmp1380;
	wire signed [31:0] w_sys_tmp1381;
	wire signed [31:0] w_sys_tmp1454;
	wire               w_sys_tmp1455;
	wire               w_sys_tmp1456;
	wire signed [31:0] w_sys_tmp1457;
	wire signed [31:0] w_sys_tmp1458;
	wire               w_sys_tmp1459;
	wire               w_sys_tmp1460;
	wire signed [31:0] w_sys_tmp1461;
	wire signed [31:0] w_sys_tmp1464;
	wire signed [31:0] w_sys_tmp1465;
	wire signed [31:0] w_sys_tmp1466;
	wire        [31:0] w_sys_tmp1467;
	wire signed [31:0] w_sys_tmp1468;
	wire signed [31:0] w_sys_tmp1469;
	wire signed [31:0] w_sys_tmp1471;
	wire signed [31:0] w_sys_tmp1472;
	wire signed [31:0] w_sys_tmp1533;
	wire               w_sys_tmp1534;
	wire               w_sys_tmp1535;
	wire signed [31:0] w_sys_tmp1536;
	wire signed [31:0] w_sys_tmp1538;
	wire signed [31:0] w_sys_tmp1539;
	wire signed [31:0] w_sys_tmp1541;
	wire signed [31:0] w_sys_tmp1542;
	wire signed [31:0] w_sys_tmp1543;
	wire        [31:0] w_sys_tmp1544;
	wire signed [31:0] w_sys_tmp1545;
	wire signed [31:0] w_sys_tmp1546;
	wire signed [31:0] w_sys_tmp1548;
	wire signed [31:0] w_sys_tmp1549;
	wire signed [31:0] w_sys_tmp1622;
	wire               w_sys_tmp1623;
	wire               w_sys_tmp1624;
	wire signed [31:0] w_sys_tmp1625;
	wire signed [31:0] w_sys_tmp1627;
	wire signed [31:0] w_sys_tmp1628;
	wire signed [31:0] w_sys_tmp1630;
	wire signed [31:0] w_sys_tmp1631;
	wire signed [31:0] w_sys_tmp1632;
	wire        [31:0] w_sys_tmp1633;
	wire signed [31:0] w_sys_tmp1634;
	wire signed [31:0] w_sys_tmp1635;
	wire signed [31:0] w_sys_tmp1637;
	wire signed [31:0] w_sys_tmp1638;
	wire signed [31:0] w_sys_tmp1711;
	wire               w_sys_tmp1712;
	wire               w_sys_tmp1713;
	wire signed [31:0] w_sys_tmp1714;
	wire signed [31:0] w_sys_tmp1716;
	wire signed [31:0] w_sys_tmp1717;
	wire signed [31:0] w_sys_tmp1719;
	wire signed [31:0] w_sys_tmp1720;
	wire signed [31:0] w_sys_tmp1721;
	wire        [31:0] w_sys_tmp1722;
	wire signed [31:0] w_sys_tmp1723;
	wire signed [31:0] w_sys_tmp1724;
	wire signed [31:0] w_sys_tmp1726;
	wire signed [31:0] w_sys_tmp1727;
	wire signed [31:0] w_sys_tmp1800;
	wire               w_sys_tmp1801;
	wire               w_sys_tmp1802;
	wire signed [31:0] w_sys_tmp1803;
	wire signed [31:0] w_sys_tmp1805;
	wire signed [31:0] w_sys_tmp1806;
	wire signed [31:0] w_sys_tmp1808;
	wire signed [31:0] w_sys_tmp1809;
	wire signed [31:0] w_sys_tmp1810;
	wire        [31:0] w_sys_tmp1811;
	wire signed [31:0] w_sys_tmp1812;
	wire signed [31:0] w_sys_tmp1813;
	wire signed [31:0] w_sys_tmp1815;
	wire signed [31:0] w_sys_tmp1816;
	wire signed [31:0] w_sys_tmp1889;
	wire               w_sys_tmp1890;
	wire               w_sys_tmp1891;
	wire signed [31:0] w_sys_tmp1892;
	wire signed [31:0] w_sys_tmp1894;
	wire signed [31:0] w_sys_tmp1895;
	wire signed [31:0] w_sys_tmp1897;
	wire signed [31:0] w_sys_tmp1898;
	wire signed [31:0] w_sys_tmp1899;
	wire        [31:0] w_sys_tmp1900;
	wire signed [31:0] w_sys_tmp1901;
	wire signed [31:0] w_sys_tmp1902;
	wire signed [31:0] w_sys_tmp1904;
	wire signed [31:0] w_sys_tmp1905;
	wire signed [31:0] w_sys_tmp1978;
	wire               w_sys_tmp1979;
	wire               w_sys_tmp1980;
	wire signed [31:0] w_sys_tmp1981;
	wire signed [31:0] w_sys_tmp1983;
	wire signed [31:0] w_sys_tmp1984;
	wire signed [31:0] w_sys_tmp1986;
	wire signed [31:0] w_sys_tmp1987;
	wire signed [31:0] w_sys_tmp1988;
	wire        [31:0] w_sys_tmp1989;
	wire signed [31:0] w_sys_tmp1990;
	wire signed [31:0] w_sys_tmp1991;
	wire signed [31:0] w_sys_tmp1993;
	wire signed [31:0] w_sys_tmp1994;
	wire signed [31:0] w_sys_tmp2067;
	wire               w_sys_tmp2068;
	wire               w_sys_tmp2069;
	wire signed [31:0] w_sys_tmp2070;
	wire signed [31:0] w_sys_tmp2072;
	wire signed [31:0] w_sys_tmp2073;
	wire signed [31:0] w_sys_tmp2075;
	wire signed [31:0] w_sys_tmp2076;
	wire signed [31:0] w_sys_tmp2077;
	wire        [31:0] w_sys_tmp2078;
	wire signed [31:0] w_sys_tmp2079;
	wire signed [31:0] w_sys_tmp2080;
	wire signed [31:0] w_sys_tmp2082;
	wire signed [31:0] w_sys_tmp2083;
	wire signed [31:0] w_sys_tmp2156;
	wire               w_sys_tmp2157;
	wire               w_sys_tmp2158;
	wire signed [31:0] w_sys_tmp2159;
	wire signed [31:0] w_sys_tmp2160;
	wire               w_sys_tmp2161;
	wire               w_sys_tmp2162;
	wire signed [31:0] w_sys_tmp2163;
	wire signed [31:0] w_sys_tmp2166;
	wire signed [31:0] w_sys_tmp2167;
	wire signed [31:0] w_sys_tmp2168;
	wire        [31:0] w_sys_tmp2169;
	wire signed [31:0] w_sys_tmp2170;
	wire signed [31:0] w_sys_tmp2171;
	wire signed [31:0] w_sys_tmp2173;
	wire signed [31:0] w_sys_tmp2174;
	wire signed [31:0] w_sys_tmp2235;
	wire               w_sys_tmp2236;
	wire               w_sys_tmp2237;
	wire signed [31:0] w_sys_tmp2238;
	wire signed [31:0] w_sys_tmp2240;
	wire signed [31:0] w_sys_tmp2241;
	wire signed [31:0] w_sys_tmp2243;
	wire signed [31:0] w_sys_tmp2244;
	wire signed [31:0] w_sys_tmp2245;
	wire        [31:0] w_sys_tmp2246;
	wire signed [31:0] w_sys_tmp2247;
	wire signed [31:0] w_sys_tmp2248;
	wire signed [31:0] w_sys_tmp2250;
	wire signed [31:0] w_sys_tmp2251;
	wire signed [31:0] w_sys_tmp2324;
	wire               w_sys_tmp2325;
	wire               w_sys_tmp2326;
	wire signed [31:0] w_sys_tmp2327;
	wire signed [31:0] w_sys_tmp2329;
	wire signed [31:0] w_sys_tmp2330;
	wire signed [31:0] w_sys_tmp2332;
	wire signed [31:0] w_sys_tmp2333;
	wire signed [31:0] w_sys_tmp2334;
	wire        [31:0] w_sys_tmp2335;
	wire signed [31:0] w_sys_tmp2336;
	wire signed [31:0] w_sys_tmp2337;
	wire signed [31:0] w_sys_tmp2339;
	wire signed [31:0] w_sys_tmp2340;
	wire signed [31:0] w_sys_tmp2413;
	wire               w_sys_tmp2414;
	wire               w_sys_tmp2415;
	wire signed [31:0] w_sys_tmp2416;
	wire signed [31:0] w_sys_tmp2418;
	wire signed [31:0] w_sys_tmp2419;
	wire signed [31:0] w_sys_tmp2421;
	wire signed [31:0] w_sys_tmp2422;
	wire signed [31:0] w_sys_tmp2423;
	wire        [31:0] w_sys_tmp2424;
	wire signed [31:0] w_sys_tmp2425;
	wire signed [31:0] w_sys_tmp2426;
	wire signed [31:0] w_sys_tmp2428;
	wire signed [31:0] w_sys_tmp2429;
	wire signed [31:0] w_sys_tmp2502;
	wire               w_sys_tmp2503;
	wire               w_sys_tmp2504;
	wire signed [31:0] w_sys_tmp2505;
	wire signed [31:0] w_sys_tmp2507;
	wire signed [31:0] w_sys_tmp2508;
	wire signed [31:0] w_sys_tmp2510;
	wire signed [31:0] w_sys_tmp2511;
	wire signed [31:0] w_sys_tmp2512;
	wire        [31:0] w_sys_tmp2513;
	wire signed [31:0] w_sys_tmp2514;
	wire signed [31:0] w_sys_tmp2515;
	wire signed [31:0] w_sys_tmp2517;
	wire signed [31:0] w_sys_tmp2518;
	wire signed [31:0] w_sys_tmp2591;
	wire               w_sys_tmp2592;
	wire               w_sys_tmp2593;
	wire signed [31:0] w_sys_tmp2594;
	wire signed [31:0] w_sys_tmp2596;
	wire signed [31:0] w_sys_tmp2597;
	wire signed [31:0] w_sys_tmp2599;
	wire signed [31:0] w_sys_tmp2600;
	wire signed [31:0] w_sys_tmp2601;
	wire        [31:0] w_sys_tmp2602;
	wire signed [31:0] w_sys_tmp2603;
	wire signed [31:0] w_sys_tmp2604;
	wire signed [31:0] w_sys_tmp2606;
	wire signed [31:0] w_sys_tmp2607;
	wire signed [31:0] w_sys_tmp2680;
	wire               w_sys_tmp2681;
	wire               w_sys_tmp2682;
	wire signed [31:0] w_sys_tmp2683;
	wire signed [31:0] w_sys_tmp2685;
	wire signed [31:0] w_sys_tmp2686;
	wire signed [31:0] w_sys_tmp2688;
	wire signed [31:0] w_sys_tmp2689;
	wire signed [31:0] w_sys_tmp2690;
	wire        [31:0] w_sys_tmp2691;
	wire signed [31:0] w_sys_tmp2692;
	wire signed [31:0] w_sys_tmp2693;
	wire signed [31:0] w_sys_tmp2695;
	wire signed [31:0] w_sys_tmp2696;
	wire signed [31:0] w_sys_tmp2769;
	wire               w_sys_tmp2770;
	wire               w_sys_tmp2771;
	wire signed [31:0] w_sys_tmp2772;
	wire signed [31:0] w_sys_tmp2774;
	wire signed [31:0] w_sys_tmp2775;
	wire signed [31:0] w_sys_tmp2777;
	wire signed [31:0] w_sys_tmp2778;
	wire signed [31:0] w_sys_tmp2779;
	wire        [31:0] w_sys_tmp2780;
	wire signed [31:0] w_sys_tmp2781;
	wire signed [31:0] w_sys_tmp2782;
	wire signed [31:0] w_sys_tmp2784;
	wire signed [31:0] w_sys_tmp2785;
	wire               w_sys_tmp2858;
	wire               w_sys_tmp2859;
	wire signed [31:0] w_sys_tmp2860;
	wire signed [31:0] w_sys_tmp2861;
	wire               w_sys_tmp2862;
	wire               w_sys_tmp2863;
	wire signed [31:0] w_sys_tmp2864;
	wire signed [31:0] w_sys_tmp2867;
	wire signed [31:0] w_sys_tmp2868;
	wire        [31:0] w_sys_tmp2869;
	wire signed [31:0] w_sys_tmp2870;
	wire signed [31:0] w_sys_tmp2871;
	wire signed [31:0] w_sys_tmp2873;
	wire signed [31:0] w_sys_tmp2874;
	wire        [31:0] w_sys_tmp2875;
	wire signed [31:0] w_sys_tmp2876;
	wire signed [31:0] w_sys_tmp2877;
	wire signed [31:0] w_sys_tmp2879;
	wire signed [31:0] w_sys_tmp2880;
	wire        [31:0] w_sys_tmp2897;
	wire        [31:0] w_sys_tmp2908;
	wire        [31:0] w_sys_tmp2919;
	wire        [31:0] w_sys_tmp2930;
	wire        [31:0] w_sys_tmp2941;
	wire signed [31:0] w_sys_tmp2944;
	wire signed [31:0] w_sys_tmp2945;
	wire               w_sys_tmp2946;
	wire               w_sys_tmp2947;
	wire signed [31:0] w_sys_tmp2948;
	wire signed [31:0] w_sys_tmp2951;
	wire signed [31:0] w_sys_tmp2952;
	wire        [31:0] w_sys_tmp2953;
	wire signed [31:0] w_sys_tmp2954;
	wire signed [31:0] w_sys_tmp2955;
	wire signed [31:0] w_sys_tmp2957;
	wire signed [31:0] w_sys_tmp2958;
	wire        [31:0] w_sys_tmp2959;
	wire signed [31:0] w_sys_tmp2960;
	wire signed [31:0] w_sys_tmp2961;
	wire signed [31:0] w_sys_tmp2963;
	wire signed [31:0] w_sys_tmp2964;
	wire        [31:0] w_sys_tmp2981;
	wire        [31:0] w_sys_tmp2992;
	wire        [31:0] w_sys_tmp3003;
	wire        [31:0] w_sys_tmp3014;
	wire        [31:0] w_sys_tmp3025;
	wire signed [31:0] w_sys_tmp3028;
	wire signed [31:0] w_sys_tmp3029;
	wire               w_sys_tmp3030;
	wire               w_sys_tmp3031;
	wire signed [31:0] w_sys_tmp3032;
	wire signed [31:0] w_sys_tmp3035;
	wire signed [31:0] w_sys_tmp3036;
	wire        [31:0] w_sys_tmp3037;
	wire signed [31:0] w_sys_tmp3038;
	wire signed [31:0] w_sys_tmp3039;
	wire signed [31:0] w_sys_tmp3041;
	wire signed [31:0] w_sys_tmp3042;
	wire        [31:0] w_sys_tmp3043;
	wire signed [31:0] w_sys_tmp3044;
	wire signed [31:0] w_sys_tmp3045;
	wire signed [31:0] w_sys_tmp3047;
	wire signed [31:0] w_sys_tmp3048;
	wire        [31:0] w_sys_tmp3065;
	wire        [31:0] w_sys_tmp3076;
	wire        [31:0] w_sys_tmp3087;
	wire        [31:0] w_sys_tmp3098;
	wire        [31:0] w_sys_tmp3109;
	wire signed [31:0] w_sys_tmp3112;
	wire signed [31:0] w_sys_tmp3113;
	wire               w_sys_tmp3114;
	wire               w_sys_tmp3115;
	wire signed [31:0] w_sys_tmp3116;
	wire signed [31:0] w_sys_tmp3119;
	wire signed [31:0] w_sys_tmp3120;
	wire        [31:0] w_sys_tmp3121;
	wire signed [31:0] w_sys_tmp3122;
	wire signed [31:0] w_sys_tmp3123;
	wire signed [31:0] w_sys_tmp3125;
	wire signed [31:0] w_sys_tmp3126;
	wire        [31:0] w_sys_tmp3127;
	wire signed [31:0] w_sys_tmp3128;
	wire signed [31:0] w_sys_tmp3129;
	wire signed [31:0] w_sys_tmp3131;
	wire signed [31:0] w_sys_tmp3132;
	wire        [31:0] w_sys_tmp3149;
	wire        [31:0] w_sys_tmp3160;
	wire        [31:0] w_sys_tmp3171;
	wire        [31:0] w_sys_tmp3182;
	wire        [31:0] w_sys_tmp3193;
	wire signed [31:0] w_sys_tmp3196;
	wire               w_sys_tmp3197;
	wire               w_sys_tmp3198;
	wire signed [31:0] w_sys_tmp3199;
	wire signed [31:0] w_sys_tmp3202;
	wire signed [31:0] w_sys_tmp3203;
	wire signed [31:0] w_sys_tmp3204;
	wire signed [31:0] w_sys_tmp3205;
	wire        [31:0] w_sys_tmp3206;
	wire signed [31:0] w_sys_tmp3207;
	wire signed [31:0] w_sys_tmp3208;
	wire signed [31:0] w_sys_tmp3212;
	wire signed [31:0] w_sys_tmp3213;
	wire signed [31:0] w_sys_tmp3215;
	wire        [31:0] w_sys_tmp3216;
	wire signed [31:0] w_sys_tmp3217;
	wire signed [31:0] w_sys_tmp3218;
	wire signed [31:0] w_sys_tmp3222;
	wire signed [31:0] w_sys_tmp3223;
	wire signed [31:0] w_sys_tmp3225;
	wire signed [31:0] w_sys_tmp3226;
	wire signed [31:0] w_sys_tmp3227;
	wire signed [31:0] w_sys_tmp3231;
	wire signed [31:0] w_sys_tmp3232;
	wire signed [31:0] w_sys_tmp3234;
	wire signed [31:0] w_sys_tmp3236;
	wire signed [31:0] w_sys_tmp3237;
	wire signed [31:0] w_sys_tmp3241;
	wire signed [31:0] w_sys_tmp3242;
	wire signed [31:0] w_sys_tmp3244;
	wire signed [31:0] w_sys_tmp3245;
	wire signed [31:0] w_sys_tmp3246;
	wire signed [31:0] w_sys_tmp3250;
	wire signed [31:0] w_sys_tmp3251;
	wire signed [31:0] w_sys_tmp3253;
	wire        [31:0] w_sys_tmp3254;
	wire signed [31:0] w_sys_tmp3255;
	wire signed [31:0] w_sys_tmp3256;
	wire signed [31:0] w_sys_tmp3259;
	wire signed [31:0] w_sys_tmp3260;
	wire signed [31:0] w_sys_tmp3261;
	wire signed [31:0] w_sys_tmp3262;
	wire signed [31:0] w_sys_tmp3263;
	wire signed [31:0] w_sys_tmp3264;
	wire signed [31:0] w_sys_tmp3265;
	wire signed [31:0] w_sys_tmp3266;
	wire signed [31:0] w_sys_tmp3267;
	wire signed [31:0] w_sys_tmp3268;
	wire signed [31:0] w_sys_tmp3269;
	wire signed [31:0] w_sys_tmp3270;
	wire signed [31:0] w_sys_tmp3697;
	wire               w_sys_tmp3698;
	wire               w_sys_tmp3699;
	wire signed [31:0] w_sys_tmp3700;
	wire signed [31:0] w_sys_tmp3703;
	wire signed [31:0] w_sys_tmp3704;
	wire signed [31:0] w_sys_tmp3705;
	wire signed [31:0] w_sys_tmp3706;
	wire        [31:0] w_sys_tmp3707;
	wire signed [31:0] w_sys_tmp3708;
	wire signed [31:0] w_sys_tmp3709;
	wire signed [31:0] w_sys_tmp3713;
	wire signed [31:0] w_sys_tmp3714;
	wire signed [31:0] w_sys_tmp3716;
	wire        [31:0] w_sys_tmp3717;
	wire signed [31:0] w_sys_tmp3718;
	wire signed [31:0] w_sys_tmp3719;
	wire signed [31:0] w_sys_tmp3723;
	wire signed [31:0] w_sys_tmp3724;
	wire signed [31:0] w_sys_tmp3726;
	wire signed [31:0] w_sys_tmp3727;
	wire signed [31:0] w_sys_tmp3728;
	wire signed [31:0] w_sys_tmp3732;
	wire signed [31:0] w_sys_tmp3733;
	wire signed [31:0] w_sys_tmp3735;
	wire signed [31:0] w_sys_tmp3737;
	wire signed [31:0] w_sys_tmp3738;
	wire signed [31:0] w_sys_tmp3742;
	wire signed [31:0] w_sys_tmp3743;
	wire signed [31:0] w_sys_tmp3745;
	wire signed [31:0] w_sys_tmp3746;
	wire signed [31:0] w_sys_tmp3747;
	wire signed [31:0] w_sys_tmp3751;
	wire signed [31:0] w_sys_tmp3752;
	wire signed [31:0] w_sys_tmp3754;
	wire        [31:0] w_sys_tmp3755;
	wire signed [31:0] w_sys_tmp3756;
	wire signed [31:0] w_sys_tmp3757;
	wire signed [31:0] w_sys_tmp3760;
	wire signed [31:0] w_sys_tmp3761;
	wire signed [31:0] w_sys_tmp3762;
	wire signed [31:0] w_sys_tmp3763;
	wire signed [31:0] w_sys_tmp3764;
	wire signed [31:0] w_sys_tmp3765;
	wire signed [31:0] w_sys_tmp3766;
	wire signed [31:0] w_sys_tmp3767;
	wire signed [31:0] w_sys_tmp3768;
	wire signed [31:0] w_sys_tmp3769;
	wire signed [31:0] w_sys_tmp3770;
	wire signed [31:0] w_sys_tmp3771;
	wire signed [31:0] w_sys_tmp4198;
	wire               w_sys_tmp4199;
	wire               w_sys_tmp4200;
	wire signed [31:0] w_sys_tmp4201;
	wire signed [31:0] w_sys_tmp4204;
	wire signed [31:0] w_sys_tmp4205;
	wire signed [31:0] w_sys_tmp4206;
	wire signed [31:0] w_sys_tmp4207;
	wire        [31:0] w_sys_tmp4208;
	wire signed [31:0] w_sys_tmp4209;
	wire signed [31:0] w_sys_tmp4210;
	wire signed [31:0] w_sys_tmp4214;
	wire signed [31:0] w_sys_tmp4215;
	wire signed [31:0] w_sys_tmp4217;
	wire        [31:0] w_sys_tmp4218;
	wire signed [31:0] w_sys_tmp4219;
	wire signed [31:0] w_sys_tmp4220;
	wire signed [31:0] w_sys_tmp4224;
	wire signed [31:0] w_sys_tmp4225;
	wire signed [31:0] w_sys_tmp4227;
	wire signed [31:0] w_sys_tmp4228;
	wire signed [31:0] w_sys_tmp4229;
	wire signed [31:0] w_sys_tmp4233;
	wire signed [31:0] w_sys_tmp4234;
	wire signed [31:0] w_sys_tmp4236;
	wire signed [31:0] w_sys_tmp4238;
	wire signed [31:0] w_sys_tmp4239;
	wire signed [31:0] w_sys_tmp4243;
	wire signed [31:0] w_sys_tmp4244;
	wire signed [31:0] w_sys_tmp4246;
	wire signed [31:0] w_sys_tmp4247;
	wire signed [31:0] w_sys_tmp4248;
	wire signed [31:0] w_sys_tmp4252;
	wire signed [31:0] w_sys_tmp4253;
	wire signed [31:0] w_sys_tmp4255;
	wire        [31:0] w_sys_tmp4256;
	wire signed [31:0] w_sys_tmp4257;
	wire signed [31:0] w_sys_tmp4258;
	wire signed [31:0] w_sys_tmp4261;
	wire signed [31:0] w_sys_tmp4262;
	wire signed [31:0] w_sys_tmp4263;
	wire signed [31:0] w_sys_tmp4264;
	wire signed [31:0] w_sys_tmp4265;
	wire signed [31:0] w_sys_tmp4266;
	wire signed [31:0] w_sys_tmp4267;
	wire signed [31:0] w_sys_tmp4268;
	wire signed [31:0] w_sys_tmp4269;
	wire signed [31:0] w_sys_tmp4270;
	wire signed [31:0] w_sys_tmp4271;
	wire signed [31:0] w_sys_tmp4272;
	wire signed [31:0] w_sys_tmp4699;
	wire               w_sys_tmp4700;
	wire               w_sys_tmp4701;
	wire signed [31:0] w_sys_tmp4702;
	wire signed [31:0] w_sys_tmp4705;
	wire signed [31:0] w_sys_tmp4706;
	wire signed [31:0] w_sys_tmp4707;
	wire signed [31:0] w_sys_tmp4708;
	wire        [31:0] w_sys_tmp4709;
	wire signed [31:0] w_sys_tmp4710;
	wire signed [31:0] w_sys_tmp4711;
	wire signed [31:0] w_sys_tmp4715;
	wire signed [31:0] w_sys_tmp4716;
	wire signed [31:0] w_sys_tmp4718;
	wire        [31:0] w_sys_tmp4719;
	wire signed [31:0] w_sys_tmp4720;
	wire signed [31:0] w_sys_tmp4721;
	wire signed [31:0] w_sys_tmp4725;
	wire signed [31:0] w_sys_tmp4726;
	wire signed [31:0] w_sys_tmp4728;
	wire signed [31:0] w_sys_tmp4729;
	wire signed [31:0] w_sys_tmp4730;
	wire signed [31:0] w_sys_tmp4734;
	wire signed [31:0] w_sys_tmp4735;
	wire signed [31:0] w_sys_tmp4737;
	wire signed [31:0] w_sys_tmp4739;
	wire signed [31:0] w_sys_tmp4740;
	wire signed [31:0] w_sys_tmp4744;
	wire signed [31:0] w_sys_tmp4745;
	wire signed [31:0] w_sys_tmp4747;
	wire signed [31:0] w_sys_tmp4748;
	wire signed [31:0] w_sys_tmp4749;
	wire signed [31:0] w_sys_tmp4753;
	wire signed [31:0] w_sys_tmp4754;
	wire signed [31:0] w_sys_tmp4756;
	wire        [31:0] w_sys_tmp4757;
	wire signed [31:0] w_sys_tmp4758;
	wire signed [31:0] w_sys_tmp4759;
	wire signed [31:0] w_sys_tmp4762;
	wire signed [31:0] w_sys_tmp4763;
	wire signed [31:0] w_sys_tmp4764;
	wire signed [31:0] w_sys_tmp4765;
	wire signed [31:0] w_sys_tmp4766;
	wire signed [31:0] w_sys_tmp4767;
	wire signed [31:0] w_sys_tmp4768;
	wire signed [31:0] w_sys_tmp4769;
	wire signed [31:0] w_sys_tmp4770;
	wire signed [31:0] w_sys_tmp4771;
	wire signed [31:0] w_sys_tmp4772;
	wire signed [31:0] w_sys_tmp4773;
	wire signed [31:0] w_sys_tmp5200;
	wire               w_sys_tmp5201;
	wire               w_sys_tmp5202;
	wire signed [31:0] w_sys_tmp5203;
	wire signed [31:0] w_sys_tmp5206;
	wire signed [31:0] w_sys_tmp5207;
	wire signed [31:0] w_sys_tmp5208;
	wire signed [31:0] w_sys_tmp5209;
	wire        [31:0] w_sys_tmp5210;
	wire signed [31:0] w_sys_tmp5211;
	wire signed [31:0] w_sys_tmp5212;
	wire signed [31:0] w_sys_tmp5216;
	wire signed [31:0] w_sys_tmp5217;
	wire signed [31:0] w_sys_tmp5219;
	wire        [31:0] w_sys_tmp5220;
	wire signed [31:0] w_sys_tmp5221;
	wire signed [31:0] w_sys_tmp5222;
	wire signed [31:0] w_sys_tmp5226;
	wire signed [31:0] w_sys_tmp5227;
	wire signed [31:0] w_sys_tmp5229;
	wire signed [31:0] w_sys_tmp5230;
	wire signed [31:0] w_sys_tmp5231;
	wire signed [31:0] w_sys_tmp5235;
	wire signed [31:0] w_sys_tmp5236;
	wire signed [31:0] w_sys_tmp5238;
	wire signed [31:0] w_sys_tmp5240;
	wire signed [31:0] w_sys_tmp5241;
	wire signed [31:0] w_sys_tmp5245;
	wire signed [31:0] w_sys_tmp5246;
	wire signed [31:0] w_sys_tmp5248;
	wire signed [31:0] w_sys_tmp5249;
	wire signed [31:0] w_sys_tmp5250;
	wire signed [31:0] w_sys_tmp5254;
	wire signed [31:0] w_sys_tmp5255;
	wire signed [31:0] w_sys_tmp5257;
	wire        [31:0] w_sys_tmp5258;
	wire signed [31:0] w_sys_tmp5259;
	wire signed [31:0] w_sys_tmp5260;
	wire signed [31:0] w_sys_tmp5263;
	wire signed [31:0] w_sys_tmp5264;
	wire signed [31:0] w_sys_tmp5265;
	wire signed [31:0] w_sys_tmp5266;
	wire signed [31:0] w_sys_tmp5267;
	wire signed [31:0] w_sys_tmp5268;
	wire signed [31:0] w_sys_tmp5269;
	wire signed [31:0] w_sys_tmp5270;
	wire signed [31:0] w_sys_tmp5271;
	wire signed [31:0] w_sys_tmp5272;
	wire signed [31:0] w_sys_tmp5273;
	wire signed [31:0] w_sys_tmp5274;
	wire signed [31:0] w_sys_tmp5701;
	wire               w_sys_tmp5702;
	wire               w_sys_tmp5703;
	wire signed [31:0] w_sys_tmp5704;
	wire signed [31:0] w_sys_tmp5707;
	wire signed [31:0] w_sys_tmp5708;
	wire signed [31:0] w_sys_tmp5709;
	wire signed [31:0] w_sys_tmp5710;
	wire        [31:0] w_sys_tmp5711;
	wire signed [31:0] w_sys_tmp5712;
	wire signed [31:0] w_sys_tmp5713;
	wire signed [31:0] w_sys_tmp5717;
	wire signed [31:0] w_sys_tmp5718;
	wire signed [31:0] w_sys_tmp5720;
	wire        [31:0] w_sys_tmp5721;
	wire signed [31:0] w_sys_tmp5722;
	wire signed [31:0] w_sys_tmp5723;
	wire signed [31:0] w_sys_tmp5727;
	wire signed [31:0] w_sys_tmp5728;
	wire signed [31:0] w_sys_tmp5730;
	wire signed [31:0] w_sys_tmp5731;
	wire signed [31:0] w_sys_tmp5732;
	wire signed [31:0] w_sys_tmp5736;
	wire signed [31:0] w_sys_tmp5737;
	wire signed [31:0] w_sys_tmp5739;
	wire signed [31:0] w_sys_tmp5741;
	wire signed [31:0] w_sys_tmp5742;
	wire signed [31:0] w_sys_tmp5746;
	wire signed [31:0] w_sys_tmp5747;
	wire signed [31:0] w_sys_tmp5749;
	wire signed [31:0] w_sys_tmp5750;
	wire signed [31:0] w_sys_tmp5751;
	wire signed [31:0] w_sys_tmp5755;
	wire signed [31:0] w_sys_tmp5756;
	wire signed [31:0] w_sys_tmp5758;
	wire        [31:0] w_sys_tmp5759;
	wire signed [31:0] w_sys_tmp5760;
	wire signed [31:0] w_sys_tmp5761;
	wire signed [31:0] w_sys_tmp5764;
	wire signed [31:0] w_sys_tmp5765;
	wire signed [31:0] w_sys_tmp5766;
	wire signed [31:0] w_sys_tmp5767;
	wire signed [31:0] w_sys_tmp5768;
	wire signed [31:0] w_sys_tmp5769;
	wire signed [31:0] w_sys_tmp5770;
	wire signed [31:0] w_sys_tmp5771;
	wire signed [31:0] w_sys_tmp5772;
	wire signed [31:0] w_sys_tmp5773;
	wire signed [31:0] w_sys_tmp5774;
	wire signed [31:0] w_sys_tmp5775;
	wire signed [31:0] w_sys_tmp6202;
	wire               w_sys_tmp6203;
	wire               w_sys_tmp6204;
	wire signed [31:0] w_sys_tmp6205;
	wire signed [31:0] w_sys_tmp6208;
	wire signed [31:0] w_sys_tmp6209;
	wire signed [31:0] w_sys_tmp6210;
	wire signed [31:0] w_sys_tmp6211;
	wire        [31:0] w_sys_tmp6212;
	wire signed [31:0] w_sys_tmp6213;
	wire signed [31:0] w_sys_tmp6214;
	wire signed [31:0] w_sys_tmp6218;
	wire signed [31:0] w_sys_tmp6219;
	wire signed [31:0] w_sys_tmp6221;
	wire        [31:0] w_sys_tmp6222;
	wire signed [31:0] w_sys_tmp6223;
	wire signed [31:0] w_sys_tmp6224;
	wire signed [31:0] w_sys_tmp6228;
	wire signed [31:0] w_sys_tmp6229;
	wire signed [31:0] w_sys_tmp6231;
	wire signed [31:0] w_sys_tmp6232;
	wire signed [31:0] w_sys_tmp6233;
	wire signed [31:0] w_sys_tmp6237;
	wire signed [31:0] w_sys_tmp6238;
	wire signed [31:0] w_sys_tmp6240;
	wire signed [31:0] w_sys_tmp6242;
	wire signed [31:0] w_sys_tmp6243;
	wire signed [31:0] w_sys_tmp6247;
	wire signed [31:0] w_sys_tmp6248;
	wire signed [31:0] w_sys_tmp6250;
	wire signed [31:0] w_sys_tmp6251;
	wire signed [31:0] w_sys_tmp6252;
	wire signed [31:0] w_sys_tmp6256;
	wire signed [31:0] w_sys_tmp6257;
	wire signed [31:0] w_sys_tmp6259;
	wire        [31:0] w_sys_tmp6260;
	wire signed [31:0] w_sys_tmp6261;
	wire signed [31:0] w_sys_tmp6262;
	wire signed [31:0] w_sys_tmp6265;
	wire signed [31:0] w_sys_tmp6266;
	wire signed [31:0] w_sys_tmp6267;
	wire signed [31:0] w_sys_tmp6268;
	wire signed [31:0] w_sys_tmp6269;
	wire signed [31:0] w_sys_tmp6270;
	wire signed [31:0] w_sys_tmp6271;
	wire signed [31:0] w_sys_tmp6272;
	wire signed [31:0] w_sys_tmp6273;
	wire signed [31:0] w_sys_tmp6274;
	wire signed [31:0] w_sys_tmp6275;
	wire signed [31:0] w_sys_tmp6276;
	wire signed [31:0] w_sys_tmp6703;
	wire               w_sys_tmp6704;
	wire               w_sys_tmp6705;
	wire signed [31:0] w_sys_tmp6706;
	wire signed [31:0] w_sys_tmp6709;
	wire signed [31:0] w_sys_tmp6710;
	wire signed [31:0] w_sys_tmp6711;
	wire signed [31:0] w_sys_tmp6712;
	wire        [31:0] w_sys_tmp6713;
	wire signed [31:0] w_sys_tmp6714;
	wire signed [31:0] w_sys_tmp6715;
	wire signed [31:0] w_sys_tmp6719;
	wire signed [31:0] w_sys_tmp6720;
	wire signed [31:0] w_sys_tmp6722;
	wire        [31:0] w_sys_tmp6723;
	wire signed [31:0] w_sys_tmp6724;
	wire signed [31:0] w_sys_tmp6725;
	wire signed [31:0] w_sys_tmp6729;
	wire signed [31:0] w_sys_tmp6730;
	wire signed [31:0] w_sys_tmp6732;
	wire signed [31:0] w_sys_tmp6733;
	wire signed [31:0] w_sys_tmp6734;
	wire signed [31:0] w_sys_tmp6738;
	wire signed [31:0] w_sys_tmp6739;
	wire signed [31:0] w_sys_tmp6741;
	wire signed [31:0] w_sys_tmp6743;
	wire signed [31:0] w_sys_tmp6744;
	wire signed [31:0] w_sys_tmp6748;
	wire signed [31:0] w_sys_tmp6749;
	wire signed [31:0] w_sys_tmp6751;
	wire signed [31:0] w_sys_tmp6752;
	wire signed [31:0] w_sys_tmp6753;
	wire signed [31:0] w_sys_tmp6757;
	wire signed [31:0] w_sys_tmp6758;
	wire signed [31:0] w_sys_tmp6760;
	wire        [31:0] w_sys_tmp6761;
	wire signed [31:0] w_sys_tmp6762;
	wire signed [31:0] w_sys_tmp6763;
	wire signed [31:0] w_sys_tmp6766;
	wire signed [31:0] w_sys_tmp6767;
	wire signed [31:0] w_sys_tmp6768;
	wire signed [31:0] w_sys_tmp6769;
	wire signed [31:0] w_sys_tmp6770;
	wire signed [31:0] w_sys_tmp6771;
	wire signed [31:0] w_sys_tmp6772;
	wire signed [31:0] w_sys_tmp6773;
	wire signed [31:0] w_sys_tmp6774;
	wire signed [31:0] w_sys_tmp6775;
	wire signed [31:0] w_sys_tmp6776;
	wire signed [31:0] w_sys_tmp6777;
	wire signed [31:0] w_sys_tmp7192;
	wire               w_sys_tmp7193;
	wire               w_sys_tmp7194;
	wire signed [31:0] w_sys_tmp7195;
	wire signed [31:0] w_sys_tmp7196;
	wire signed [31:0] w_sys_tmp7197;
	wire               w_sys_tmp7198;
	wire               w_sys_tmp7199;
	wire signed [31:0] w_sys_tmp7200;
	wire signed [31:0] w_sys_tmp7203;
	wire signed [31:0] w_sys_tmp7204;
	wire signed [31:0] w_sys_tmp7205;
	wire        [31:0] w_sys_tmp7206;
	wire signed [31:0] w_sys_tmp7207;
	wire signed [31:0] w_sys_tmp7208;
	wire signed [31:0] w_sys_tmp7210;
	wire signed [31:0] w_sys_tmp7211;
	wire signed [31:0] w_sys_tmp7272;
	wire               w_sys_tmp7273;
	wire               w_sys_tmp7274;
	wire signed [31:0] w_sys_tmp7275;
	wire signed [31:0] w_sys_tmp7277;
	wire signed [31:0] w_sys_tmp7278;
	wire signed [31:0] w_sys_tmp7280;
	wire signed [31:0] w_sys_tmp7281;
	wire signed [31:0] w_sys_tmp7282;
	wire        [31:0] w_sys_tmp7283;
	wire signed [31:0] w_sys_tmp7284;
	wire signed [31:0] w_sys_tmp7285;
	wire signed [31:0] w_sys_tmp7287;
	wire signed [31:0] w_sys_tmp7288;
	wire signed [31:0] w_sys_tmp7289;
	wire signed [31:0] w_sys_tmp7368;
	wire               w_sys_tmp7369;
	wire               w_sys_tmp7370;
	wire signed [31:0] w_sys_tmp7371;
	wire signed [31:0] w_sys_tmp7373;
	wire signed [31:0] w_sys_tmp7374;
	wire signed [31:0] w_sys_tmp7376;
	wire signed [31:0] w_sys_tmp7377;
	wire signed [31:0] w_sys_tmp7378;
	wire        [31:0] w_sys_tmp7379;
	wire signed [31:0] w_sys_tmp7380;
	wire signed [31:0] w_sys_tmp7381;
	wire signed [31:0] w_sys_tmp7383;
	wire signed [31:0] w_sys_tmp7384;
	wire signed [31:0] w_sys_tmp7385;
	wire signed [31:0] w_sys_tmp7464;
	wire               w_sys_tmp7465;
	wire               w_sys_tmp7466;
	wire signed [31:0] w_sys_tmp7467;
	wire signed [31:0] w_sys_tmp7469;
	wire signed [31:0] w_sys_tmp7470;
	wire signed [31:0] w_sys_tmp7472;
	wire signed [31:0] w_sys_tmp7473;
	wire signed [31:0] w_sys_tmp7474;
	wire        [31:0] w_sys_tmp7475;
	wire signed [31:0] w_sys_tmp7476;
	wire signed [31:0] w_sys_tmp7477;
	wire signed [31:0] w_sys_tmp7479;
	wire signed [31:0] w_sys_tmp7480;
	wire signed [31:0] w_sys_tmp7481;
	wire signed [31:0] w_sys_tmp7560;
	wire               w_sys_tmp7561;
	wire               w_sys_tmp7562;
	wire signed [31:0] w_sys_tmp7563;
	wire signed [31:0] w_sys_tmp7565;
	wire signed [31:0] w_sys_tmp7566;
	wire signed [31:0] w_sys_tmp7568;
	wire signed [31:0] w_sys_tmp7569;
	wire signed [31:0] w_sys_tmp7570;
	wire        [31:0] w_sys_tmp7571;
	wire signed [31:0] w_sys_tmp7572;
	wire signed [31:0] w_sys_tmp7573;
	wire signed [31:0] w_sys_tmp7575;
	wire signed [31:0] w_sys_tmp7576;
	wire signed [31:0] w_sys_tmp7577;
	wire signed [31:0] w_sys_tmp7656;
	wire               w_sys_tmp7657;
	wire               w_sys_tmp7658;
	wire signed [31:0] w_sys_tmp7659;
	wire signed [31:0] w_sys_tmp7661;
	wire signed [31:0] w_sys_tmp7662;
	wire signed [31:0] w_sys_tmp7664;
	wire signed [31:0] w_sys_tmp7665;
	wire signed [31:0] w_sys_tmp7666;
	wire        [31:0] w_sys_tmp7667;
	wire signed [31:0] w_sys_tmp7668;
	wire signed [31:0] w_sys_tmp7669;
	wire signed [31:0] w_sys_tmp7671;
	wire signed [31:0] w_sys_tmp7672;
	wire signed [31:0] w_sys_tmp7673;
	wire signed [31:0] w_sys_tmp7752;
	wire               w_sys_tmp7753;
	wire               w_sys_tmp7754;
	wire signed [31:0] w_sys_tmp7755;
	wire signed [31:0] w_sys_tmp7757;
	wire signed [31:0] w_sys_tmp7758;
	wire signed [31:0] w_sys_tmp7760;
	wire signed [31:0] w_sys_tmp7761;
	wire signed [31:0] w_sys_tmp7762;
	wire        [31:0] w_sys_tmp7763;
	wire signed [31:0] w_sys_tmp7764;
	wire signed [31:0] w_sys_tmp7765;
	wire signed [31:0] w_sys_tmp7767;
	wire signed [31:0] w_sys_tmp7768;
	wire signed [31:0] w_sys_tmp7769;
	wire signed [31:0] w_sys_tmp7848;
	wire               w_sys_tmp7849;
	wire               w_sys_tmp7850;
	wire signed [31:0] w_sys_tmp7851;
	wire signed [31:0] w_sys_tmp7853;
	wire signed [31:0] w_sys_tmp7854;
	wire signed [31:0] w_sys_tmp7856;
	wire signed [31:0] w_sys_tmp7857;
	wire signed [31:0] w_sys_tmp7858;
	wire        [31:0] w_sys_tmp7859;
	wire signed [31:0] w_sys_tmp7860;
	wire signed [31:0] w_sys_tmp7861;
	wire signed [31:0] w_sys_tmp7863;
	wire signed [31:0] w_sys_tmp7864;
	wire signed [31:0] w_sys_tmp7865;
	wire signed [31:0] w_sys_tmp7944;
	wire               w_sys_tmp7945;
	wire               w_sys_tmp7946;
	wire signed [31:0] w_sys_tmp7947;
	wire signed [31:0] w_sys_tmp7948;
	wire signed [31:0] w_sys_tmp7949;
	wire               w_sys_tmp7950;
	wire               w_sys_tmp7951;
	wire signed [31:0] w_sys_tmp7952;
	wire signed [31:0] w_sys_tmp7955;
	wire signed [31:0] w_sys_tmp7956;
	wire signed [31:0] w_sys_tmp7957;
	wire        [31:0] w_sys_tmp7958;
	wire signed [31:0] w_sys_tmp7959;
	wire signed [31:0] w_sys_tmp7960;
	wire signed [31:0] w_sys_tmp7962;
	wire signed [31:0] w_sys_tmp7963;
	wire signed [31:0] w_sys_tmp8024;
	wire               w_sys_tmp8025;
	wire               w_sys_tmp8026;
	wire signed [31:0] w_sys_tmp8027;
	wire signed [31:0] w_sys_tmp8029;
	wire signed [31:0] w_sys_tmp8030;
	wire signed [31:0] w_sys_tmp8032;
	wire signed [31:0] w_sys_tmp8033;
	wire signed [31:0] w_sys_tmp8034;
	wire        [31:0] w_sys_tmp8035;
	wire signed [31:0] w_sys_tmp8036;
	wire signed [31:0] w_sys_tmp8037;
	wire signed [31:0] w_sys_tmp8039;
	wire signed [31:0] w_sys_tmp8040;
	wire signed [31:0] w_sys_tmp8041;
	wire signed [31:0] w_sys_tmp8120;
	wire               w_sys_tmp8121;
	wire               w_sys_tmp8122;
	wire signed [31:0] w_sys_tmp8123;
	wire signed [31:0] w_sys_tmp8125;
	wire signed [31:0] w_sys_tmp8126;
	wire signed [31:0] w_sys_tmp8128;
	wire signed [31:0] w_sys_tmp8129;
	wire signed [31:0] w_sys_tmp8130;
	wire        [31:0] w_sys_tmp8131;
	wire signed [31:0] w_sys_tmp8132;
	wire signed [31:0] w_sys_tmp8133;
	wire signed [31:0] w_sys_tmp8135;
	wire signed [31:0] w_sys_tmp8136;
	wire signed [31:0] w_sys_tmp8137;
	wire signed [31:0] w_sys_tmp8216;
	wire               w_sys_tmp8217;
	wire               w_sys_tmp8218;
	wire signed [31:0] w_sys_tmp8219;
	wire signed [31:0] w_sys_tmp8221;
	wire signed [31:0] w_sys_tmp8222;
	wire signed [31:0] w_sys_tmp8224;
	wire signed [31:0] w_sys_tmp8225;
	wire signed [31:0] w_sys_tmp8226;
	wire        [31:0] w_sys_tmp8227;
	wire signed [31:0] w_sys_tmp8228;
	wire signed [31:0] w_sys_tmp8229;
	wire signed [31:0] w_sys_tmp8231;
	wire signed [31:0] w_sys_tmp8232;
	wire signed [31:0] w_sys_tmp8233;
	wire signed [31:0] w_sys_tmp8312;
	wire               w_sys_tmp8313;
	wire               w_sys_tmp8314;
	wire signed [31:0] w_sys_tmp8315;
	wire signed [31:0] w_sys_tmp8317;
	wire signed [31:0] w_sys_tmp8318;
	wire signed [31:0] w_sys_tmp8320;
	wire signed [31:0] w_sys_tmp8321;
	wire signed [31:0] w_sys_tmp8322;
	wire        [31:0] w_sys_tmp8323;
	wire signed [31:0] w_sys_tmp8324;
	wire signed [31:0] w_sys_tmp8325;
	wire signed [31:0] w_sys_tmp8327;
	wire signed [31:0] w_sys_tmp8328;
	wire signed [31:0] w_sys_tmp8329;
	wire signed [31:0] w_sys_tmp8408;
	wire               w_sys_tmp8409;
	wire               w_sys_tmp8410;
	wire signed [31:0] w_sys_tmp8411;
	wire signed [31:0] w_sys_tmp8413;
	wire signed [31:0] w_sys_tmp8414;
	wire signed [31:0] w_sys_tmp8416;
	wire signed [31:0] w_sys_tmp8417;
	wire signed [31:0] w_sys_tmp8418;
	wire        [31:0] w_sys_tmp8419;
	wire signed [31:0] w_sys_tmp8420;
	wire signed [31:0] w_sys_tmp8421;
	wire signed [31:0] w_sys_tmp8423;
	wire signed [31:0] w_sys_tmp8424;
	wire signed [31:0] w_sys_tmp8425;
	wire signed [31:0] w_sys_tmp8504;
	wire               w_sys_tmp8505;
	wire               w_sys_tmp8506;
	wire signed [31:0] w_sys_tmp8507;
	wire signed [31:0] w_sys_tmp8509;
	wire signed [31:0] w_sys_tmp8510;
	wire signed [31:0] w_sys_tmp8512;
	wire signed [31:0] w_sys_tmp8513;
	wire signed [31:0] w_sys_tmp8514;
	wire        [31:0] w_sys_tmp8515;
	wire signed [31:0] w_sys_tmp8516;
	wire signed [31:0] w_sys_tmp8517;
	wire signed [31:0] w_sys_tmp8519;
	wire signed [31:0] w_sys_tmp8520;
	wire signed [31:0] w_sys_tmp8521;
	wire signed [31:0] w_sys_tmp8600;
	wire               w_sys_tmp8601;
	wire               w_sys_tmp8602;
	wire signed [31:0] w_sys_tmp8603;
	wire signed [31:0] w_sys_tmp8605;
	wire signed [31:0] w_sys_tmp8606;
	wire signed [31:0] w_sys_tmp8608;
	wire signed [31:0] w_sys_tmp8609;
	wire signed [31:0] w_sys_tmp8610;
	wire        [31:0] w_sys_tmp8611;
	wire signed [31:0] w_sys_tmp8612;
	wire signed [31:0] w_sys_tmp8613;
	wire signed [31:0] w_sys_tmp8615;
	wire signed [31:0] w_sys_tmp8616;
	wire signed [31:0] w_sys_tmp8617;
	wire signed [31:0] w_sys_tmp8696;
	wire               w_sys_tmp8697;
	wire               w_sys_tmp8698;
	wire signed [31:0] w_sys_tmp8699;
	wire signed [31:0] w_sys_tmp8700;
	wire signed [31:0] w_sys_tmp8701;
	wire               w_sys_tmp8702;
	wire               w_sys_tmp8703;
	wire signed [31:0] w_sys_tmp8704;
	wire signed [31:0] w_sys_tmp8707;
	wire signed [31:0] w_sys_tmp8708;
	wire signed [31:0] w_sys_tmp8709;
	wire        [31:0] w_sys_tmp8710;
	wire signed [31:0] w_sys_tmp8711;
	wire signed [31:0] w_sys_tmp8712;
	wire signed [31:0] w_sys_tmp8714;
	wire signed [31:0] w_sys_tmp8715;
	wire signed [31:0] w_sys_tmp8776;
	wire               w_sys_tmp8777;
	wire               w_sys_tmp8778;
	wire signed [31:0] w_sys_tmp8779;
	wire signed [31:0] w_sys_tmp8781;
	wire signed [31:0] w_sys_tmp8782;
	wire signed [31:0] w_sys_tmp8784;
	wire signed [31:0] w_sys_tmp8785;
	wire signed [31:0] w_sys_tmp8786;
	wire        [31:0] w_sys_tmp8787;
	wire signed [31:0] w_sys_tmp8788;
	wire signed [31:0] w_sys_tmp8789;
	wire signed [31:0] w_sys_tmp8791;
	wire signed [31:0] w_sys_tmp8792;
	wire signed [31:0] w_sys_tmp8793;
	wire signed [31:0] w_sys_tmp8872;
	wire               w_sys_tmp8873;
	wire               w_sys_tmp8874;
	wire signed [31:0] w_sys_tmp8875;
	wire signed [31:0] w_sys_tmp8877;
	wire signed [31:0] w_sys_tmp8878;
	wire signed [31:0] w_sys_tmp8880;
	wire signed [31:0] w_sys_tmp8881;
	wire signed [31:0] w_sys_tmp8882;
	wire        [31:0] w_sys_tmp8883;
	wire signed [31:0] w_sys_tmp8884;
	wire signed [31:0] w_sys_tmp8885;
	wire signed [31:0] w_sys_tmp8887;
	wire signed [31:0] w_sys_tmp8888;
	wire signed [31:0] w_sys_tmp8889;
	wire signed [31:0] w_sys_tmp8968;
	wire               w_sys_tmp8969;
	wire               w_sys_tmp8970;
	wire signed [31:0] w_sys_tmp8971;
	wire signed [31:0] w_sys_tmp8973;
	wire signed [31:0] w_sys_tmp8974;
	wire signed [31:0] w_sys_tmp8976;
	wire signed [31:0] w_sys_tmp8977;
	wire signed [31:0] w_sys_tmp8978;
	wire        [31:0] w_sys_tmp8979;
	wire signed [31:0] w_sys_tmp8980;
	wire signed [31:0] w_sys_tmp8981;
	wire signed [31:0] w_sys_tmp8983;
	wire signed [31:0] w_sys_tmp8984;
	wire signed [31:0] w_sys_tmp8985;
	wire signed [31:0] w_sys_tmp9064;
	wire               w_sys_tmp9065;
	wire               w_sys_tmp9066;
	wire signed [31:0] w_sys_tmp9067;
	wire signed [31:0] w_sys_tmp9069;
	wire signed [31:0] w_sys_tmp9070;
	wire signed [31:0] w_sys_tmp9072;
	wire signed [31:0] w_sys_tmp9073;
	wire signed [31:0] w_sys_tmp9074;
	wire        [31:0] w_sys_tmp9075;
	wire signed [31:0] w_sys_tmp9076;
	wire signed [31:0] w_sys_tmp9077;
	wire signed [31:0] w_sys_tmp9079;
	wire signed [31:0] w_sys_tmp9080;
	wire signed [31:0] w_sys_tmp9081;
	wire signed [31:0] w_sys_tmp9160;
	wire               w_sys_tmp9161;
	wire               w_sys_tmp9162;
	wire signed [31:0] w_sys_tmp9163;
	wire signed [31:0] w_sys_tmp9165;
	wire signed [31:0] w_sys_tmp9166;
	wire signed [31:0] w_sys_tmp9168;
	wire signed [31:0] w_sys_tmp9169;
	wire signed [31:0] w_sys_tmp9170;
	wire        [31:0] w_sys_tmp9171;
	wire signed [31:0] w_sys_tmp9172;
	wire signed [31:0] w_sys_tmp9173;
	wire signed [31:0] w_sys_tmp9175;
	wire signed [31:0] w_sys_tmp9176;
	wire signed [31:0] w_sys_tmp9177;
	wire signed [31:0] w_sys_tmp9256;
	wire               w_sys_tmp9257;
	wire               w_sys_tmp9258;
	wire signed [31:0] w_sys_tmp9259;
	wire signed [31:0] w_sys_tmp9261;
	wire signed [31:0] w_sys_tmp9262;
	wire signed [31:0] w_sys_tmp9264;
	wire signed [31:0] w_sys_tmp9265;
	wire signed [31:0] w_sys_tmp9266;
	wire        [31:0] w_sys_tmp9267;
	wire signed [31:0] w_sys_tmp9268;
	wire signed [31:0] w_sys_tmp9269;
	wire signed [31:0] w_sys_tmp9271;
	wire signed [31:0] w_sys_tmp9272;
	wire signed [31:0] w_sys_tmp9273;
	wire signed [31:0] w_sys_tmp9352;
	wire               w_sys_tmp9353;
	wire               w_sys_tmp9354;
	wire signed [31:0] w_sys_tmp9355;
	wire signed [31:0] w_sys_tmp9357;
	wire signed [31:0] w_sys_tmp9358;
	wire signed [31:0] w_sys_tmp9360;
	wire signed [31:0] w_sys_tmp9361;
	wire signed [31:0] w_sys_tmp9362;
	wire        [31:0] w_sys_tmp9363;
	wire signed [31:0] w_sys_tmp9364;
	wire signed [31:0] w_sys_tmp9365;
	wire signed [31:0] w_sys_tmp9367;
	wire signed [31:0] w_sys_tmp9368;
	wire signed [31:0] w_sys_tmp9369;
	wire signed [31:0] w_sys_tmp9448;
	wire               w_sys_tmp9449;
	wire               w_sys_tmp9450;
	wire signed [31:0] w_sys_tmp9451;
	wire signed [31:0] w_sys_tmp9452;
	wire signed [31:0] w_sys_tmp9453;
	wire               w_sys_tmp9454;
	wire               w_sys_tmp9455;
	wire signed [31:0] w_sys_tmp9456;
	wire signed [31:0] w_sys_tmp9459;
	wire signed [31:0] w_sys_tmp9460;
	wire signed [31:0] w_sys_tmp9461;
	wire        [31:0] w_sys_tmp9462;
	wire signed [31:0] w_sys_tmp9463;
	wire signed [31:0] w_sys_tmp9464;
	wire signed [31:0] w_sys_tmp9466;
	wire signed [31:0] w_sys_tmp9467;
	wire signed [31:0] w_sys_tmp9528;
	wire               w_sys_tmp9529;
	wire               w_sys_tmp9530;
	wire signed [31:0] w_sys_tmp9531;
	wire signed [31:0] w_sys_tmp9533;
	wire signed [31:0] w_sys_tmp9534;
	wire signed [31:0] w_sys_tmp9536;
	wire signed [31:0] w_sys_tmp9537;
	wire signed [31:0] w_sys_tmp9538;
	wire        [31:0] w_sys_tmp9539;
	wire signed [31:0] w_sys_tmp9540;
	wire signed [31:0] w_sys_tmp9541;
	wire signed [31:0] w_sys_tmp9543;
	wire signed [31:0] w_sys_tmp9544;
	wire signed [31:0] w_sys_tmp9545;
	wire signed [31:0] w_sys_tmp9624;
	wire               w_sys_tmp9625;
	wire               w_sys_tmp9626;
	wire signed [31:0] w_sys_tmp9627;
	wire signed [31:0] w_sys_tmp9629;
	wire signed [31:0] w_sys_tmp9630;
	wire signed [31:0] w_sys_tmp9632;
	wire signed [31:0] w_sys_tmp9633;
	wire signed [31:0] w_sys_tmp9634;
	wire        [31:0] w_sys_tmp9635;
	wire signed [31:0] w_sys_tmp9636;
	wire signed [31:0] w_sys_tmp9637;
	wire signed [31:0] w_sys_tmp9639;
	wire signed [31:0] w_sys_tmp9640;
	wire signed [31:0] w_sys_tmp9641;
	wire signed [31:0] w_sys_tmp9720;
	wire               w_sys_tmp9721;
	wire               w_sys_tmp9722;
	wire signed [31:0] w_sys_tmp9723;
	wire signed [31:0] w_sys_tmp9725;
	wire signed [31:0] w_sys_tmp9726;
	wire signed [31:0] w_sys_tmp9728;
	wire signed [31:0] w_sys_tmp9729;
	wire signed [31:0] w_sys_tmp9730;
	wire        [31:0] w_sys_tmp9731;
	wire signed [31:0] w_sys_tmp9732;
	wire signed [31:0] w_sys_tmp9733;
	wire signed [31:0] w_sys_tmp9735;
	wire signed [31:0] w_sys_tmp9736;
	wire signed [31:0] w_sys_tmp9737;
	wire signed [31:0] w_sys_tmp9816;
	wire               w_sys_tmp9817;
	wire               w_sys_tmp9818;
	wire signed [31:0] w_sys_tmp9819;
	wire signed [31:0] w_sys_tmp9821;
	wire signed [31:0] w_sys_tmp9822;
	wire signed [31:0] w_sys_tmp9824;
	wire signed [31:0] w_sys_tmp9825;
	wire signed [31:0] w_sys_tmp9826;
	wire        [31:0] w_sys_tmp9827;
	wire signed [31:0] w_sys_tmp9828;
	wire signed [31:0] w_sys_tmp9829;
	wire signed [31:0] w_sys_tmp9831;
	wire signed [31:0] w_sys_tmp9832;
	wire signed [31:0] w_sys_tmp9833;
	wire signed [31:0] w_sys_tmp9912;
	wire               w_sys_tmp9913;
	wire               w_sys_tmp9914;
	wire signed [31:0] w_sys_tmp9915;
	wire signed [31:0] w_sys_tmp9917;
	wire signed [31:0] w_sys_tmp9918;
	wire signed [31:0] w_sys_tmp9920;
	wire signed [31:0] w_sys_tmp9921;
	wire signed [31:0] w_sys_tmp9922;
	wire        [31:0] w_sys_tmp9923;
	wire signed [31:0] w_sys_tmp9924;
	wire signed [31:0] w_sys_tmp9925;
	wire signed [31:0] w_sys_tmp9927;
	wire signed [31:0] w_sys_tmp9928;
	wire signed [31:0] w_sys_tmp9929;
	wire signed [31:0] w_sys_tmp10008;
	wire               w_sys_tmp10009;
	wire               w_sys_tmp10010;
	wire signed [31:0] w_sys_tmp10011;
	wire signed [31:0] w_sys_tmp10013;
	wire signed [31:0] w_sys_tmp10014;
	wire signed [31:0] w_sys_tmp10016;
	wire signed [31:0] w_sys_tmp10017;
	wire signed [31:0] w_sys_tmp10018;
	wire        [31:0] w_sys_tmp10019;
	wire signed [31:0] w_sys_tmp10020;
	wire signed [31:0] w_sys_tmp10021;
	wire signed [31:0] w_sys_tmp10023;
	wire signed [31:0] w_sys_tmp10024;
	wire signed [31:0] w_sys_tmp10025;
	wire signed [31:0] w_sys_tmp10104;
	wire               w_sys_tmp10105;
	wire               w_sys_tmp10106;
	wire signed [31:0] w_sys_tmp10107;
	wire signed [31:0] w_sys_tmp10109;
	wire signed [31:0] w_sys_tmp10110;
	wire signed [31:0] w_sys_tmp10112;
	wire signed [31:0] w_sys_tmp10113;
	wire signed [31:0] w_sys_tmp10114;
	wire        [31:0] w_sys_tmp10115;
	wire signed [31:0] w_sys_tmp10116;
	wire signed [31:0] w_sys_tmp10117;
	wire signed [31:0] w_sys_tmp10119;
	wire signed [31:0] w_sys_tmp10120;
	wire signed [31:0] w_sys_tmp10121;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 6'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 6'h1);
	assign w_fld_u_0_addr_0 = 15'sh0;
	assign w_fld_u_0_datain_0 = 32'h0;
	assign w_fld_u_0_r_w_0 = 1'h0;
	assign w_fld_u_0_ce_0 = w_sys_ce;
	assign w_fld_u_0_ce_1 = w_sys_ce;
	assign w_sub19_u_addr = ( (|r_sys_processing_methodID) ? r_sub19_u_addr : 12'sh0 ) ;
	assign w_sub19_u_datain = ( (|r_sys_processing_methodID) ? r_sub19_u_datain : 32'h0 ) ;
	assign w_sub19_u_r_w = ( (|r_sys_processing_methodID) ? r_sub19_u_r_w : 1'h0 ) ;
	assign w_sub19_result_addr = ( (|r_sys_processing_methodID) ? r_sub19_result_addr : 12'sh0 ) ;
	assign w_sub19_result_datain = ( (|r_sys_processing_methodID) ? r_sub19_result_datain : 32'h0 ) ;
	assign w_sub19_result_r_w = ( (|r_sys_processing_methodID) ? r_sub19_result_r_w : 1'h0 ) ;
	assign w_sub12_u_addr = ( (|r_sys_processing_methodID) ? r_sub12_u_addr : 12'sh0 ) ;
	assign w_sub12_u_datain = ( (|r_sys_processing_methodID) ? r_sub12_u_datain : 32'h0 ) ;
	assign w_sub12_u_r_w = ( (|r_sys_processing_methodID) ? r_sub12_u_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 12'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub11_u_addr = ( (|r_sys_processing_methodID) ? r_sub11_u_addr : 12'sh0 ) ;
	assign w_sub11_u_datain = ( (|r_sys_processing_methodID) ? r_sub11_u_datain : 32'h0 ) ;
	assign w_sub11_u_r_w = ( (|r_sys_processing_methodID) ? r_sub11_u_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 12'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_u_addr = ( (|r_sys_processing_methodID) ? r_sub14_u_addr : 12'sh0 ) ;
	assign w_sub14_u_datain = ( (|r_sys_processing_methodID) ? r_sub14_u_datain : 32'h0 ) ;
	assign w_sub14_u_r_w = ( (|r_sys_processing_methodID) ? r_sub14_u_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 12'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub13_u_addr = ( (|r_sys_processing_methodID) ? r_sub13_u_addr : 12'sh0 ) ;
	assign w_sub13_u_datain = ( (|r_sys_processing_methodID) ? r_sub13_u_datain : 32'h0 ) ;
	assign w_sub13_u_r_w = ( (|r_sys_processing_methodID) ? r_sub13_u_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 12'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub16_u_addr = ( (|r_sys_processing_methodID) ? r_sub16_u_addr : 12'sh0 ) ;
	assign w_sub16_u_datain = ( (|r_sys_processing_methodID) ? r_sub16_u_datain : 32'h0 ) ;
	assign w_sub16_u_r_w = ( (|r_sys_processing_methodID) ? r_sub16_u_r_w : 1'h0 ) ;
	assign w_sub16_result_addr = ( (|r_sys_processing_methodID) ? r_sub16_result_addr : 12'sh0 ) ;
	assign w_sub16_result_datain = ( (|r_sys_processing_methodID) ? r_sub16_result_datain : 32'h0 ) ;
	assign w_sub16_result_r_w = ( (|r_sys_processing_methodID) ? r_sub16_result_r_w : 1'h0 ) ;
	assign w_sub15_u_addr = ( (|r_sys_processing_methodID) ? r_sub15_u_addr : 12'sh0 ) ;
	assign w_sub15_u_datain = ( (|r_sys_processing_methodID) ? r_sub15_u_datain : 32'h0 ) ;
	assign w_sub15_u_r_w = ( (|r_sys_processing_methodID) ? r_sub15_u_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 12'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub18_u_addr = ( (|r_sys_processing_methodID) ? r_sub18_u_addr : 12'sh0 ) ;
	assign w_sub18_u_datain = ( (|r_sys_processing_methodID) ? r_sub18_u_datain : 32'h0 ) ;
	assign w_sub18_u_r_w = ( (|r_sys_processing_methodID) ? r_sub18_u_r_w : 1'h0 ) ;
	assign w_sub18_result_addr = ( (|r_sys_processing_methodID) ? r_sub18_result_addr : 12'sh0 ) ;
	assign w_sub18_result_datain = ( (|r_sys_processing_methodID) ? r_sub18_result_datain : 32'h0 ) ;
	assign w_sub18_result_r_w = ( (|r_sys_processing_methodID) ? r_sub18_result_r_w : 1'h0 ) ;
	assign w_sub17_u_addr = ( (|r_sys_processing_methodID) ? r_sub17_u_addr : 12'sh0 ) ;
	assign w_sub17_u_datain = ( (|r_sys_processing_methodID) ? r_sub17_u_datain : 32'h0 ) ;
	assign w_sub17_u_r_w = ( (|r_sys_processing_methodID) ? r_sub17_u_r_w : 1'h0 ) ;
	assign w_sub17_result_addr = ( (|r_sys_processing_methodID) ? r_sub17_result_addr : 12'sh0 ) ;
	assign w_sub17_result_datain = ( (|r_sys_processing_methodID) ? r_sub17_result_datain : 32'h0 ) ;
	assign w_sub17_result_r_w = ( (|r_sys_processing_methodID) ? r_sub17_result_r_w : 1'h0 ) ;
	assign w_sub20_u_addr = ( (|r_sys_processing_methodID) ? r_sub20_u_addr : 12'sh0 ) ;
	assign w_sub20_u_datain = ( (|r_sys_processing_methodID) ? r_sub20_u_datain : 32'h0 ) ;
	assign w_sub20_u_r_w = ( (|r_sys_processing_methodID) ? r_sub20_u_r_w : 1'h0 ) ;
	assign w_sub20_result_addr = ( (|r_sys_processing_methodID) ? r_sub20_result_addr : 12'sh0 ) ;
	assign w_sub20_result_datain = ( (|r_sys_processing_methodID) ? r_sub20_result_datain : 32'h0 ) ;
	assign w_sub20_result_r_w = ( (|r_sys_processing_methodID) ? r_sub20_result_r_w : 1'h0 ) ;
	assign w_sub21_u_addr = ( (|r_sys_processing_methodID) ? r_sub21_u_addr : 12'sh0 ) ;
	assign w_sub21_u_datain = ( (|r_sys_processing_methodID) ? r_sub21_u_datain : 32'h0 ) ;
	assign w_sub21_u_r_w = ( (|r_sys_processing_methodID) ? r_sub21_u_r_w : 1'h0 ) ;
	assign w_sub21_result_addr = ( (|r_sys_processing_methodID) ? r_sub21_result_addr : 12'sh0 ) ;
	assign w_sub21_result_datain = ( (|r_sys_processing_methodID) ? r_sub21_result_datain : 32'h0 ) ;
	assign w_sub21_result_r_w = ( (|r_sys_processing_methodID) ? r_sub21_result_r_w : 1'h0 ) ;
	assign w_sub28_u_addr = ( (|r_sys_processing_methodID) ? r_sub28_u_addr : 12'sh0 ) ;
	assign w_sub28_u_datain = ( (|r_sys_processing_methodID) ? r_sub28_u_datain : 32'h0 ) ;
	assign w_sub28_u_r_w = ( (|r_sys_processing_methodID) ? r_sub28_u_r_w : 1'h0 ) ;
	assign w_sub28_result_addr = ( (|r_sys_processing_methodID) ? r_sub28_result_addr : 12'sh0 ) ;
	assign w_sub28_result_datain = ( (|r_sys_processing_methodID) ? r_sub28_result_datain : 32'h0 ) ;
	assign w_sub28_result_r_w = ( (|r_sys_processing_methodID) ? r_sub28_result_r_w : 1'h0 ) ;
	assign w_sub29_u_addr = ( (|r_sys_processing_methodID) ? r_sub29_u_addr : 12'sh0 ) ;
	assign w_sub29_u_datain = ( (|r_sys_processing_methodID) ? r_sub29_u_datain : 32'h0 ) ;
	assign w_sub29_u_r_w = ( (|r_sys_processing_methodID) ? r_sub29_u_r_w : 1'h0 ) ;
	assign w_sub29_result_addr = ( (|r_sys_processing_methodID) ? r_sub29_result_addr : 12'sh0 ) ;
	assign w_sub29_result_datain = ( (|r_sys_processing_methodID) ? r_sub29_result_datain : 32'h0 ) ;
	assign w_sub29_result_r_w = ( (|r_sys_processing_methodID) ? r_sub29_result_r_w : 1'h0 ) ;
	assign w_sub26_u_addr = ( (|r_sys_processing_methodID) ? r_sub26_u_addr : 12'sh0 ) ;
	assign w_sub26_u_datain = ( (|r_sys_processing_methodID) ? r_sub26_u_datain : 32'h0 ) ;
	assign w_sub26_u_r_w = ( (|r_sys_processing_methodID) ? r_sub26_u_r_w : 1'h0 ) ;
	assign w_sub26_result_addr = ( (|r_sys_processing_methodID) ? r_sub26_result_addr : 12'sh0 ) ;
	assign w_sub26_result_datain = ( (|r_sys_processing_methodID) ? r_sub26_result_datain : 32'h0 ) ;
	assign w_sub26_result_r_w = ( (|r_sys_processing_methodID) ? r_sub26_result_r_w : 1'h0 ) ;
	assign w_sub09_u_addr = ( (|r_sys_processing_methodID) ? r_sub09_u_addr : 12'sh0 ) ;
	assign w_sub09_u_datain = ( (|r_sys_processing_methodID) ? r_sub09_u_datain : 32'h0 ) ;
	assign w_sub09_u_r_w = ( (|r_sys_processing_methodID) ? r_sub09_u_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 12'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub27_u_addr = ( (|r_sys_processing_methodID) ? r_sub27_u_addr : 12'sh0 ) ;
	assign w_sub27_u_datain = ( (|r_sys_processing_methodID) ? r_sub27_u_datain : 32'h0 ) ;
	assign w_sub27_u_r_w = ( (|r_sys_processing_methodID) ? r_sub27_u_r_w : 1'h0 ) ;
	assign w_sub27_result_addr = ( (|r_sys_processing_methodID) ? r_sub27_result_addr : 12'sh0 ) ;
	assign w_sub27_result_datain = ( (|r_sys_processing_methodID) ? r_sub27_result_datain : 32'h0 ) ;
	assign w_sub27_result_r_w = ( (|r_sys_processing_methodID) ? r_sub27_result_r_w : 1'h0 ) ;
	assign w_sub08_u_addr = ( (|r_sys_processing_methodID) ? r_sub08_u_addr : 12'sh0 ) ;
	assign w_sub08_u_datain = ( (|r_sys_processing_methodID) ? r_sub08_u_datain : 32'h0 ) ;
	assign w_sub08_u_r_w = ( (|r_sys_processing_methodID) ? r_sub08_u_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 12'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub24_u_addr = ( (|r_sys_processing_methodID) ? r_sub24_u_addr : 12'sh0 ) ;
	assign w_sub24_u_datain = ( (|r_sys_processing_methodID) ? r_sub24_u_datain : 32'h0 ) ;
	assign w_sub24_u_r_w = ( (|r_sys_processing_methodID) ? r_sub24_u_r_w : 1'h0 ) ;
	assign w_sub24_result_addr = ( (|r_sys_processing_methodID) ? r_sub24_result_addr : 12'sh0 ) ;
	assign w_sub24_result_datain = ( (|r_sys_processing_methodID) ? r_sub24_result_datain : 32'h0 ) ;
	assign w_sub24_result_r_w = ( (|r_sys_processing_methodID) ? r_sub24_result_r_w : 1'h0 ) ;
	assign w_sub25_u_addr = ( (|r_sys_processing_methodID) ? r_sub25_u_addr : 12'sh0 ) ;
	assign w_sub25_u_datain = ( (|r_sys_processing_methodID) ? r_sub25_u_datain : 32'h0 ) ;
	assign w_sub25_u_r_w = ( (|r_sys_processing_methodID) ? r_sub25_u_r_w : 1'h0 ) ;
	assign w_sub25_result_addr = ( (|r_sys_processing_methodID) ? r_sub25_result_addr : 12'sh0 ) ;
	assign w_sub25_result_datain = ( (|r_sys_processing_methodID) ? r_sub25_result_datain : 32'h0 ) ;
	assign w_sub25_result_r_w = ( (|r_sys_processing_methodID) ? r_sub25_result_r_w : 1'h0 ) ;
	assign w_sub22_u_addr = ( (|r_sys_processing_methodID) ? r_sub22_u_addr : 12'sh0 ) ;
	assign w_sub22_u_datain = ( (|r_sys_processing_methodID) ? r_sub22_u_datain : 32'h0 ) ;
	assign w_sub22_u_r_w = ( (|r_sys_processing_methodID) ? r_sub22_u_r_w : 1'h0 ) ;
	assign w_sub22_result_addr = ( (|r_sys_processing_methodID) ? r_sub22_result_addr : 12'sh0 ) ;
	assign w_sub22_result_datain = ( (|r_sys_processing_methodID) ? r_sub22_result_datain : 32'h0 ) ;
	assign w_sub22_result_r_w = ( (|r_sys_processing_methodID) ? r_sub22_result_r_w : 1'h0 ) ;
	assign w_sub23_u_addr = ( (|r_sys_processing_methodID) ? r_sub23_u_addr : 12'sh0 ) ;
	assign w_sub23_u_datain = ( (|r_sys_processing_methodID) ? r_sub23_u_datain : 32'h0 ) ;
	assign w_sub23_u_r_w = ( (|r_sys_processing_methodID) ? r_sub23_u_r_w : 1'h0 ) ;
	assign w_sub23_result_addr = ( (|r_sys_processing_methodID) ? r_sub23_result_addr : 12'sh0 ) ;
	assign w_sub23_result_datain = ( (|r_sys_processing_methodID) ? r_sub23_result_datain : 32'h0 ) ;
	assign w_sub23_result_r_w = ( (|r_sys_processing_methodID) ? r_sub23_result_r_w : 1'h0 ) ;
	assign w_sub03_u_addr = ( (|r_sys_processing_methodID) ? r_sub03_u_addr : 12'sh0 ) ;
	assign w_sub03_u_datain = ( (|r_sys_processing_methodID) ? r_sub03_u_datain : 32'h0 ) ;
	assign w_sub03_u_r_w = ( (|r_sys_processing_methodID) ? r_sub03_u_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 12'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_u_addr = ( (|r_sys_processing_methodID) ? r_sub02_u_addr : 12'sh0 ) ;
	assign w_sub02_u_datain = ( (|r_sys_processing_methodID) ? r_sub02_u_datain : 32'h0 ) ;
	assign w_sub02_u_r_w = ( (|r_sys_processing_methodID) ? r_sub02_u_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 12'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_u_addr = ( (|r_sys_processing_methodID) ? r_sub01_u_addr : 12'sh0 ) ;
	assign w_sub01_u_datain = ( (|r_sys_processing_methodID) ? r_sub01_u_datain : 32'h0 ) ;
	assign w_sub01_u_r_w = ( (|r_sys_processing_methodID) ? r_sub01_u_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 12'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_u_addr = ( (|r_sys_processing_methodID) ? r_sub00_u_addr : 12'sh0 ) ;
	assign w_sub00_u_datain = ( (|r_sys_processing_methodID) ? r_sub00_u_datain : 32'h0 ) ;
	assign w_sub00_u_r_w = ( (|r_sys_processing_methodID) ? r_sub00_u_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 12'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_u_addr = ( (|r_sys_processing_methodID) ? r_sub07_u_addr : 12'sh0 ) ;
	assign w_sub07_u_datain = ( (|r_sys_processing_methodID) ? r_sub07_u_datain : 32'h0 ) ;
	assign w_sub07_u_r_w = ( (|r_sys_processing_methodID) ? r_sub07_u_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 12'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_u_addr = ( (|r_sys_processing_methodID) ? r_sub06_u_addr : 12'sh0 ) ;
	assign w_sub06_u_datain = ( (|r_sys_processing_methodID) ? r_sub06_u_datain : 32'h0 ) ;
	assign w_sub06_u_r_w = ( (|r_sys_processing_methodID) ? r_sub06_u_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 12'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub05_u_addr = ( (|r_sys_processing_methodID) ? r_sub05_u_addr : 12'sh0 ) ;
	assign w_sub05_u_datain = ( (|r_sys_processing_methodID) ? r_sub05_u_datain : 32'h0 ) ;
	assign w_sub05_u_r_w = ( (|r_sys_processing_methodID) ? r_sub05_u_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 12'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_u_addr = ( (|r_sys_processing_methodID) ? r_sub04_u_addr : 12'sh0 ) ;
	assign w_sub04_u_datain = ( (|r_sys_processing_methodID) ? r_sub04_u_datain : 32'h0 ) ;
	assign w_sub04_u_r_w = ( (|r_sys_processing_methodID) ? r_sub04_u_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 12'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub10_u_addr = ( (|r_sys_processing_methodID) ? r_sub10_u_addr : 12'sh0 ) ;
	assign w_sub10_u_datain = ( (|r_sys_processing_methodID) ? r_sub10_u_datain : 32'h0 ) ;
	assign w_sub10_u_r_w = ( (|r_sys_processing_methodID) ? r_sub10_u_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 12'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sub31_u_addr = ( (|r_sys_processing_methodID) ? r_sub31_u_addr : 12'sh0 ) ;
	assign w_sub31_u_datain = ( (|r_sys_processing_methodID) ? r_sub31_u_datain : 32'h0 ) ;
	assign w_sub31_u_r_w = ( (|r_sys_processing_methodID) ? r_sub31_u_r_w : 1'h0 ) ;
	assign w_sub31_result_addr = ( (|r_sys_processing_methodID) ? r_sub31_result_addr : 12'sh0 ) ;
	assign w_sub31_result_datain = ( (|r_sys_processing_methodID) ? r_sub31_result_datain : 32'h0 ) ;
	assign w_sub31_result_r_w = ( (|r_sys_processing_methodID) ? r_sub31_result_r_w : 1'h0 ) ;
	assign w_sub30_u_addr = ( (|r_sys_processing_methodID) ? r_sub30_u_addr : 12'sh0 ) ;
	assign w_sub30_u_datain = ( (|r_sys_processing_methodID) ? r_sub30_u_datain : 32'h0 ) ;
	assign w_sub30_u_r_w = ( (|r_sys_processing_methodID) ? r_sub30_u_r_w : 1'h0 ) ;
	assign w_sub30_result_addr = ( (|r_sys_processing_methodID) ? r_sub30_result_addr : 12'sh0 ) ;
	assign w_sub30_result_datain = ( (|r_sys_processing_methodID) ? r_sub30_result_datain : 32'h0 ) ;
	assign w_sub30_result_r_w = ( (|r_sys_processing_methodID) ? r_sub30_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000081;
	assign w_sys_tmp3 = ( !w_sys_tmp4 );
	assign w_sys_tmp4 = (r_run_my_37 < r_run_k_33);
	assign w_sys_tmp5 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp6 = ( !w_sys_tmp7 );
	assign w_sys_tmp7 = (r_run_mx_36 < r_run_j_34);
	assign w_sys_tmp10 = (w_sys_tmp11 + r_run_k_33);
	assign w_sys_tmp11 = (r_run_j_34 * w_sys_tmp12);
	assign w_sys_tmp12 = 32'sh00000081;
	assign w_sys_tmp13 = 32'h0;
	assign w_sys_tmp14 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp51 = ( !w_sys_tmp52 );
	assign w_sys_tmp52 = (w_sys_tmp53 < r_run_k_33);
	assign w_sys_tmp53 = 32'sh00000021;
	assign w_sys_tmp54 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp55 = ( !w_sys_tmp56 );
	assign w_sys_tmp56 = (w_sys_tmp57 < r_run_j_34);
	assign w_sys_tmp57 = 32'sh00000011;
	assign w_sys_tmp60 = (w_sys_tmp61 + r_run_k_33);
	assign w_sys_tmp61 = (r_run_j_34 * w_sys_tmp62);
	assign w_sys_tmp62 = 32'sh00000081;
	assign w_sys_tmp63 = w_fld_u_0_dataout_1;
	assign w_sys_tmp64 = (w_sys_tmp65 + r_run_k_33);
	assign w_sys_tmp65 = (r_run_copy0_j_40 * w_sys_tmp62);
	assign w_sys_tmp67 = (r_run_copy0_j_40 + w_sys_intOne);
	assign w_sys_tmp68 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp129 = 32'sh00000010;
	assign w_sys_tmp130 = ( !w_sys_tmp131 );
	assign w_sys_tmp131 = (w_sys_tmp132 < r_run_j_34);
	assign w_sys_tmp132 = 32'sh00000021;
	assign w_sys_tmp134 = (r_run_j_34 - w_sys_tmp135);
	assign w_sys_tmp135 = 32'sh0000000f;
	assign w_sys_tmp137 = (w_sys_tmp138 + r_run_k_33);
	assign w_sys_tmp138 = (r_run_tmpj_39 * w_sys_tmp139);
	assign w_sys_tmp139 = 32'sh00000081;
	assign w_sys_tmp140 = w_fld_u_0_dataout_1;
	assign w_sys_tmp141 = (w_sys_tmp142 + r_run_k_33);
	assign w_sys_tmp142 = (r_run_copy0_j_41 * w_sys_tmp139);
	assign w_sys_tmp144 = (r_run_copy0_j_41 + w_sys_intOne);
	assign w_sys_tmp145 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp218 = 32'sh00000020;
	assign w_sys_tmp219 = ( !w_sys_tmp220 );
	assign w_sys_tmp220 = (w_sys_tmp221 < r_run_j_34);
	assign w_sys_tmp221 = 32'sh00000031;
	assign w_sys_tmp223 = (r_run_j_34 - w_sys_tmp224);
	assign w_sys_tmp224 = 32'sh0000001f;
	assign w_sys_tmp226 = (w_sys_tmp227 + r_run_k_33);
	assign w_sys_tmp227 = (r_run_tmpj_39 * w_sys_tmp228);
	assign w_sys_tmp228 = 32'sh00000081;
	assign w_sys_tmp229 = w_fld_u_0_dataout_1;
	assign w_sys_tmp230 = (w_sys_tmp231 + r_run_k_33);
	assign w_sys_tmp231 = (r_run_copy0_j_42 * w_sys_tmp228);
	assign w_sys_tmp233 = (r_run_copy0_j_42 + w_sys_intOne);
	assign w_sys_tmp234 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp307 = 32'sh00000030;
	assign w_sys_tmp308 = ( !w_sys_tmp309 );
	assign w_sys_tmp309 = (w_sys_tmp310 < r_run_j_34);
	assign w_sys_tmp310 = 32'sh00000041;
	assign w_sys_tmp312 = (r_run_j_34 - w_sys_tmp313);
	assign w_sys_tmp313 = 32'sh0000002f;
	assign w_sys_tmp315 = (w_sys_tmp316 + r_run_k_33);
	assign w_sys_tmp316 = (r_run_tmpj_39 * w_sys_tmp317);
	assign w_sys_tmp317 = 32'sh00000081;
	assign w_sys_tmp318 = w_fld_u_0_dataout_1;
	assign w_sys_tmp319 = (w_sys_tmp320 + r_run_k_33);
	assign w_sys_tmp320 = (r_run_copy0_j_43 * w_sys_tmp317);
	assign w_sys_tmp322 = (r_run_copy0_j_43 + w_sys_intOne);
	assign w_sys_tmp323 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp396 = 32'sh00000040;
	assign w_sys_tmp397 = ( !w_sys_tmp398 );
	assign w_sys_tmp398 = (w_sys_tmp399 < r_run_j_34);
	assign w_sys_tmp399 = 32'sh00000051;
	assign w_sys_tmp401 = (r_run_j_34 - w_sys_tmp402);
	assign w_sys_tmp402 = 32'sh0000003f;
	assign w_sys_tmp404 = (w_sys_tmp405 + r_run_k_33);
	assign w_sys_tmp405 = (r_run_tmpj_39 * w_sys_tmp406);
	assign w_sys_tmp406 = 32'sh00000081;
	assign w_sys_tmp407 = w_fld_u_0_dataout_1;
	assign w_sys_tmp408 = (w_sys_tmp409 + r_run_k_33);
	assign w_sys_tmp409 = (r_run_copy0_j_44 * w_sys_tmp406);
	assign w_sys_tmp411 = (r_run_copy0_j_44 + w_sys_intOne);
	assign w_sys_tmp412 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp485 = 32'sh00000050;
	assign w_sys_tmp486 = ( !w_sys_tmp487 );
	assign w_sys_tmp487 = (w_sys_tmp488 < r_run_j_34);
	assign w_sys_tmp488 = 32'sh00000061;
	assign w_sys_tmp490 = (r_run_j_34 - w_sys_tmp491);
	assign w_sys_tmp491 = 32'sh0000004f;
	assign w_sys_tmp493 = (w_sys_tmp494 + r_run_k_33);
	assign w_sys_tmp494 = (r_run_tmpj_39 * w_sys_tmp495);
	assign w_sys_tmp495 = 32'sh00000081;
	assign w_sys_tmp496 = w_fld_u_0_dataout_1;
	assign w_sys_tmp497 = (w_sys_tmp498 + r_run_k_33);
	assign w_sys_tmp498 = (r_run_copy0_j_45 * w_sys_tmp495);
	assign w_sys_tmp500 = (r_run_copy0_j_45 + w_sys_intOne);
	assign w_sys_tmp501 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp574 = 32'sh00000060;
	assign w_sys_tmp575 = ( !w_sys_tmp576 );
	assign w_sys_tmp576 = (w_sys_tmp577 < r_run_j_34);
	assign w_sys_tmp577 = 32'sh00000071;
	assign w_sys_tmp579 = (r_run_j_34 - w_sys_tmp580);
	assign w_sys_tmp580 = 32'sh0000005f;
	assign w_sys_tmp582 = (w_sys_tmp583 + r_run_k_33);
	assign w_sys_tmp583 = (r_run_tmpj_39 * w_sys_tmp584);
	assign w_sys_tmp584 = 32'sh00000081;
	assign w_sys_tmp585 = w_fld_u_0_dataout_1;
	assign w_sys_tmp586 = (w_sys_tmp587 + r_run_k_33);
	assign w_sys_tmp587 = (r_run_copy0_j_46 * w_sys_tmp584);
	assign w_sys_tmp589 = (r_run_copy0_j_46 + w_sys_intOne);
	assign w_sys_tmp590 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp663 = 32'sh00000070;
	assign w_sys_tmp664 = ( !w_sys_tmp665 );
	assign w_sys_tmp665 = (w_sys_tmp666 < r_run_j_34);
	assign w_sys_tmp666 = 32'sh00000081;
	assign w_sys_tmp668 = (r_run_j_34 - w_sys_tmp669);
	assign w_sys_tmp669 = 32'sh0000006f;
	assign w_sys_tmp671 = (w_sys_tmp672 + r_run_k_33);
	assign w_sys_tmp672 = (r_run_tmpj_39 * w_sys_tmp673);
	assign w_sys_tmp673 = 32'sh00000081;
	assign w_sys_tmp674 = w_fld_u_0_dataout_1;
	assign w_sys_tmp675 = (w_sys_tmp676 + r_run_k_33);
	assign w_sys_tmp676 = (r_run_copy0_j_47 * w_sys_tmp673);
	assign w_sys_tmp678 = (r_run_copy0_j_47 + w_sys_intOne);
	assign w_sys_tmp679 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp752 = 32'sh00000020;
	assign w_sys_tmp753 = ( !w_sys_tmp754 );
	assign w_sys_tmp754 = (w_sys_tmp755 < r_run_k_33);
	assign w_sys_tmp755 = 32'sh00000041;
	assign w_sys_tmp756 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp757 = ( !w_sys_tmp758 );
	assign w_sys_tmp758 = (w_sys_tmp759 < r_run_j_34);
	assign w_sys_tmp759 = 32'sh00000011;
	assign w_sys_tmp762 = (w_sys_tmp763 + r_run_k_33);
	assign w_sys_tmp763 = (r_run_j_34 * w_sys_tmp764);
	assign w_sys_tmp764 = 32'sh00000081;
	assign w_sys_tmp765 = w_fld_u_0_dataout_1;
	assign w_sys_tmp766 = (w_sys_tmp767 + r_run_k_33);
	assign w_sys_tmp767 = (r_run_copy0_j_48 * w_sys_tmp764);
	assign w_sys_tmp769 = (r_run_copy0_j_48 + w_sys_intOne);
	assign w_sys_tmp770 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp831 = 32'sh00000010;
	assign w_sys_tmp832 = ( !w_sys_tmp833 );
	assign w_sys_tmp833 = (w_sys_tmp834 < r_run_j_34);
	assign w_sys_tmp834 = 32'sh00000021;
	assign w_sys_tmp836 = (r_run_j_34 - w_sys_tmp837);
	assign w_sys_tmp837 = 32'sh0000000f;
	assign w_sys_tmp839 = (w_sys_tmp840 + r_run_k_33);
	assign w_sys_tmp840 = (r_run_tmpj_39 * w_sys_tmp841);
	assign w_sys_tmp841 = 32'sh00000081;
	assign w_sys_tmp842 = w_fld_u_0_dataout_1;
	assign w_sys_tmp843 = (w_sys_tmp844 + r_run_k_33);
	assign w_sys_tmp844 = (r_run_copy0_j_49 * w_sys_tmp841);
	assign w_sys_tmp846 = (r_run_copy0_j_49 + w_sys_intOne);
	assign w_sys_tmp847 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp920 = 32'sh00000020;
	assign w_sys_tmp921 = ( !w_sys_tmp922 );
	assign w_sys_tmp922 = (w_sys_tmp923 < r_run_j_34);
	assign w_sys_tmp923 = 32'sh00000031;
	assign w_sys_tmp925 = (r_run_j_34 - w_sys_tmp926);
	assign w_sys_tmp926 = 32'sh0000001f;
	assign w_sys_tmp928 = (w_sys_tmp929 + r_run_k_33);
	assign w_sys_tmp929 = (r_run_tmpj_39 * w_sys_tmp930);
	assign w_sys_tmp930 = 32'sh00000081;
	assign w_sys_tmp931 = w_fld_u_0_dataout_1;
	assign w_sys_tmp932 = (w_sys_tmp933 + r_run_k_33);
	assign w_sys_tmp933 = (r_run_copy0_j_50 * w_sys_tmp930);
	assign w_sys_tmp935 = (r_run_copy0_j_50 + w_sys_intOne);
	assign w_sys_tmp936 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1009 = 32'sh00000030;
	assign w_sys_tmp1010 = ( !w_sys_tmp1011 );
	assign w_sys_tmp1011 = (w_sys_tmp1012 < r_run_j_34);
	assign w_sys_tmp1012 = 32'sh00000041;
	assign w_sys_tmp1014 = (r_run_j_34 - w_sys_tmp1015);
	assign w_sys_tmp1015 = 32'sh0000002f;
	assign w_sys_tmp1017 = (w_sys_tmp1018 + r_run_k_33);
	assign w_sys_tmp1018 = (r_run_tmpj_39 * w_sys_tmp1019);
	assign w_sys_tmp1019 = 32'sh00000081;
	assign w_sys_tmp1020 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1021 = (w_sys_tmp1022 + r_run_k_33);
	assign w_sys_tmp1022 = (r_run_copy0_j_51 * w_sys_tmp1019);
	assign w_sys_tmp1024 = (r_run_copy0_j_51 + w_sys_intOne);
	assign w_sys_tmp1025 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1098 = 32'sh00000040;
	assign w_sys_tmp1099 = ( !w_sys_tmp1100 );
	assign w_sys_tmp1100 = (w_sys_tmp1101 < r_run_j_34);
	assign w_sys_tmp1101 = 32'sh00000051;
	assign w_sys_tmp1103 = (r_run_j_34 - w_sys_tmp1104);
	assign w_sys_tmp1104 = 32'sh0000003f;
	assign w_sys_tmp1106 = (w_sys_tmp1107 + r_run_k_33);
	assign w_sys_tmp1107 = (r_run_tmpj_39 * w_sys_tmp1108);
	assign w_sys_tmp1108 = 32'sh00000081;
	assign w_sys_tmp1109 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1110 = (w_sys_tmp1111 + r_run_k_33);
	assign w_sys_tmp1111 = (r_run_copy0_j_52 * w_sys_tmp1108);
	assign w_sys_tmp1113 = (r_run_copy0_j_52 + w_sys_intOne);
	assign w_sys_tmp1114 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1187 = 32'sh00000050;
	assign w_sys_tmp1188 = ( !w_sys_tmp1189 );
	assign w_sys_tmp1189 = (w_sys_tmp1190 < r_run_j_34);
	assign w_sys_tmp1190 = 32'sh00000061;
	assign w_sys_tmp1192 = (r_run_j_34 - w_sys_tmp1193);
	assign w_sys_tmp1193 = 32'sh0000004f;
	assign w_sys_tmp1195 = (w_sys_tmp1196 + r_run_k_33);
	assign w_sys_tmp1196 = (r_run_tmpj_39 * w_sys_tmp1197);
	assign w_sys_tmp1197 = 32'sh00000081;
	assign w_sys_tmp1198 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1199 = (w_sys_tmp1200 + r_run_k_33);
	assign w_sys_tmp1200 = (r_run_copy0_j_53 * w_sys_tmp1197);
	assign w_sys_tmp1202 = (r_run_copy0_j_53 + w_sys_intOne);
	assign w_sys_tmp1203 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1276 = 32'sh00000060;
	assign w_sys_tmp1277 = ( !w_sys_tmp1278 );
	assign w_sys_tmp1278 = (w_sys_tmp1279 < r_run_j_34);
	assign w_sys_tmp1279 = 32'sh00000071;
	assign w_sys_tmp1281 = (r_run_j_34 - w_sys_tmp1282);
	assign w_sys_tmp1282 = 32'sh0000005f;
	assign w_sys_tmp1284 = (w_sys_tmp1285 + r_run_k_33);
	assign w_sys_tmp1285 = (r_run_tmpj_39 * w_sys_tmp1286);
	assign w_sys_tmp1286 = 32'sh00000081;
	assign w_sys_tmp1287 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1288 = (w_sys_tmp1289 + r_run_k_33);
	assign w_sys_tmp1289 = (r_run_copy0_j_54 * w_sys_tmp1286);
	assign w_sys_tmp1291 = (r_run_copy0_j_54 + w_sys_intOne);
	assign w_sys_tmp1292 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1365 = 32'sh00000070;
	assign w_sys_tmp1366 = ( !w_sys_tmp1367 );
	assign w_sys_tmp1367 = (w_sys_tmp1368 < r_run_j_34);
	assign w_sys_tmp1368 = 32'sh00000081;
	assign w_sys_tmp1370 = (r_run_j_34 - w_sys_tmp1371);
	assign w_sys_tmp1371 = 32'sh0000006f;
	assign w_sys_tmp1373 = (w_sys_tmp1374 + r_run_k_33);
	assign w_sys_tmp1374 = (r_run_tmpj_39 * w_sys_tmp1375);
	assign w_sys_tmp1375 = 32'sh00000081;
	assign w_sys_tmp1376 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1377 = (w_sys_tmp1378 + r_run_k_33);
	assign w_sys_tmp1378 = (r_run_copy0_j_55 * w_sys_tmp1375);
	assign w_sys_tmp1380 = (r_run_copy0_j_55 + w_sys_intOne);
	assign w_sys_tmp1381 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1454 = 32'sh00000040;
	assign w_sys_tmp1455 = ( !w_sys_tmp1456 );
	assign w_sys_tmp1456 = (w_sys_tmp1457 < r_run_k_33);
	assign w_sys_tmp1457 = 32'sh00000061;
	assign w_sys_tmp1458 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp1459 = ( !w_sys_tmp1460 );
	assign w_sys_tmp1460 = (w_sys_tmp1461 < r_run_j_34);
	assign w_sys_tmp1461 = 32'sh00000011;
	assign w_sys_tmp1464 = (w_sys_tmp1465 + r_run_k_33);
	assign w_sys_tmp1465 = (r_run_j_34 * w_sys_tmp1466);
	assign w_sys_tmp1466 = 32'sh00000081;
	assign w_sys_tmp1467 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1468 = (w_sys_tmp1469 + r_run_k_33);
	assign w_sys_tmp1469 = (r_run_copy0_j_56 * w_sys_tmp1466);
	assign w_sys_tmp1471 = (r_run_copy0_j_56 + w_sys_intOne);
	assign w_sys_tmp1472 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1533 = 32'sh00000010;
	assign w_sys_tmp1534 = ( !w_sys_tmp1535 );
	assign w_sys_tmp1535 = (w_sys_tmp1536 < r_run_j_34);
	assign w_sys_tmp1536 = 32'sh00000021;
	assign w_sys_tmp1538 = (r_run_j_34 - w_sys_tmp1539);
	assign w_sys_tmp1539 = 32'sh0000000f;
	assign w_sys_tmp1541 = (w_sys_tmp1542 + r_run_k_33);
	assign w_sys_tmp1542 = (r_run_tmpj_39 * w_sys_tmp1543);
	assign w_sys_tmp1543 = 32'sh00000081;
	assign w_sys_tmp1544 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1545 = (w_sys_tmp1546 + r_run_k_33);
	assign w_sys_tmp1546 = (r_run_copy0_j_57 * w_sys_tmp1543);
	assign w_sys_tmp1548 = (r_run_copy0_j_57 + w_sys_intOne);
	assign w_sys_tmp1549 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1622 = 32'sh00000020;
	assign w_sys_tmp1623 = ( !w_sys_tmp1624 );
	assign w_sys_tmp1624 = (w_sys_tmp1625 < r_run_j_34);
	assign w_sys_tmp1625 = 32'sh00000031;
	assign w_sys_tmp1627 = (r_run_j_34 - w_sys_tmp1628);
	assign w_sys_tmp1628 = 32'sh0000001f;
	assign w_sys_tmp1630 = (w_sys_tmp1631 + r_run_k_33);
	assign w_sys_tmp1631 = (r_run_tmpj_39 * w_sys_tmp1632);
	assign w_sys_tmp1632 = 32'sh00000081;
	assign w_sys_tmp1633 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1634 = (w_sys_tmp1635 + r_run_k_33);
	assign w_sys_tmp1635 = (r_run_copy0_j_58 * w_sys_tmp1632);
	assign w_sys_tmp1637 = (r_run_copy0_j_58 + w_sys_intOne);
	assign w_sys_tmp1638 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1711 = 32'sh00000030;
	assign w_sys_tmp1712 = ( !w_sys_tmp1713 );
	assign w_sys_tmp1713 = (w_sys_tmp1714 < r_run_j_34);
	assign w_sys_tmp1714 = 32'sh00000041;
	assign w_sys_tmp1716 = (r_run_j_34 - w_sys_tmp1717);
	assign w_sys_tmp1717 = 32'sh0000002f;
	assign w_sys_tmp1719 = (w_sys_tmp1720 + r_run_k_33);
	assign w_sys_tmp1720 = (r_run_tmpj_39 * w_sys_tmp1721);
	assign w_sys_tmp1721 = 32'sh00000081;
	assign w_sys_tmp1722 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1723 = (w_sys_tmp1724 + r_run_k_33);
	assign w_sys_tmp1724 = (r_run_copy0_j_59 * w_sys_tmp1721);
	assign w_sys_tmp1726 = (r_run_copy0_j_59 + w_sys_intOne);
	assign w_sys_tmp1727 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1800 = 32'sh00000040;
	assign w_sys_tmp1801 = ( !w_sys_tmp1802 );
	assign w_sys_tmp1802 = (w_sys_tmp1803 < r_run_j_34);
	assign w_sys_tmp1803 = 32'sh00000051;
	assign w_sys_tmp1805 = (r_run_j_34 - w_sys_tmp1806);
	assign w_sys_tmp1806 = 32'sh0000003f;
	assign w_sys_tmp1808 = (w_sys_tmp1809 + r_run_k_33);
	assign w_sys_tmp1809 = (r_run_tmpj_39 * w_sys_tmp1810);
	assign w_sys_tmp1810 = 32'sh00000081;
	assign w_sys_tmp1811 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1812 = (w_sys_tmp1813 + r_run_k_33);
	assign w_sys_tmp1813 = (r_run_copy0_j_60 * w_sys_tmp1810);
	assign w_sys_tmp1815 = (r_run_copy0_j_60 + w_sys_intOne);
	assign w_sys_tmp1816 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1889 = 32'sh00000050;
	assign w_sys_tmp1890 = ( !w_sys_tmp1891 );
	assign w_sys_tmp1891 = (w_sys_tmp1892 < r_run_j_34);
	assign w_sys_tmp1892 = 32'sh00000061;
	assign w_sys_tmp1894 = (r_run_j_34 - w_sys_tmp1895);
	assign w_sys_tmp1895 = 32'sh0000004f;
	assign w_sys_tmp1897 = (w_sys_tmp1898 + r_run_k_33);
	assign w_sys_tmp1898 = (r_run_tmpj_39 * w_sys_tmp1899);
	assign w_sys_tmp1899 = 32'sh00000081;
	assign w_sys_tmp1900 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1901 = (w_sys_tmp1902 + r_run_k_33);
	assign w_sys_tmp1902 = (r_run_copy0_j_61 * w_sys_tmp1899);
	assign w_sys_tmp1904 = (r_run_copy0_j_61 + w_sys_intOne);
	assign w_sys_tmp1905 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp1978 = 32'sh00000060;
	assign w_sys_tmp1979 = ( !w_sys_tmp1980 );
	assign w_sys_tmp1980 = (w_sys_tmp1981 < r_run_j_34);
	assign w_sys_tmp1981 = 32'sh00000071;
	assign w_sys_tmp1983 = (r_run_j_34 - w_sys_tmp1984);
	assign w_sys_tmp1984 = 32'sh0000005f;
	assign w_sys_tmp1986 = (w_sys_tmp1987 + r_run_k_33);
	assign w_sys_tmp1987 = (r_run_tmpj_39 * w_sys_tmp1988);
	assign w_sys_tmp1988 = 32'sh00000081;
	assign w_sys_tmp1989 = w_fld_u_0_dataout_1;
	assign w_sys_tmp1990 = (w_sys_tmp1991 + r_run_k_33);
	assign w_sys_tmp1991 = (r_run_copy0_j_62 * w_sys_tmp1988);
	assign w_sys_tmp1993 = (r_run_copy0_j_62 + w_sys_intOne);
	assign w_sys_tmp1994 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp2067 = 32'sh00000070;
	assign w_sys_tmp2068 = ( !w_sys_tmp2069 );
	assign w_sys_tmp2069 = (w_sys_tmp2070 < r_run_j_34);
	assign w_sys_tmp2070 = 32'sh00000081;
	assign w_sys_tmp2072 = (r_run_j_34 - w_sys_tmp2073);
	assign w_sys_tmp2073 = 32'sh0000006f;
	assign w_sys_tmp2075 = (w_sys_tmp2076 + r_run_k_33);
	assign w_sys_tmp2076 = (r_run_tmpj_39 * w_sys_tmp2077);
	assign w_sys_tmp2077 = 32'sh00000081;
	assign w_sys_tmp2078 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2079 = (w_sys_tmp2080 + r_run_k_33);
	assign w_sys_tmp2080 = (r_run_copy0_j_63 * w_sys_tmp2077);
	assign w_sys_tmp2082 = (r_run_copy0_j_63 + w_sys_intOne);
	assign w_sys_tmp2083 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp2156 = 32'sh00000060;
	assign w_sys_tmp2157 = ( !w_sys_tmp2158 );
	assign w_sys_tmp2158 = (w_sys_tmp2159 < r_run_k_33);
	assign w_sys_tmp2159 = 32'sh00000081;
	assign w_sys_tmp2160 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp2161 = ( !w_sys_tmp2162 );
	assign w_sys_tmp2162 = (w_sys_tmp2163 < r_run_j_34);
	assign w_sys_tmp2163 = 32'sh00000011;
	assign w_sys_tmp2166 = (w_sys_tmp2167 + r_run_k_33);
	assign w_sys_tmp2167 = (r_run_j_34 * w_sys_tmp2168);
	assign w_sys_tmp2168 = 32'sh00000081;
	assign w_sys_tmp2169 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2170 = (w_sys_tmp2171 + r_run_k_33);
	assign w_sys_tmp2171 = (r_run_copy0_j_64 * w_sys_tmp2168);
	assign w_sys_tmp2173 = (r_run_copy0_j_64 + w_sys_intOne);
	assign w_sys_tmp2174 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp2235 = 32'sh00000010;
	assign w_sys_tmp2236 = ( !w_sys_tmp2237 );
	assign w_sys_tmp2237 = (w_sys_tmp2238 < r_run_j_34);
	assign w_sys_tmp2238 = 32'sh00000021;
	assign w_sys_tmp2240 = (r_run_j_34 - w_sys_tmp2241);
	assign w_sys_tmp2241 = 32'sh0000000f;
	assign w_sys_tmp2243 = (w_sys_tmp2244 + r_run_k_33);
	assign w_sys_tmp2244 = (r_run_tmpj_39 * w_sys_tmp2245);
	assign w_sys_tmp2245 = 32'sh00000081;
	assign w_sys_tmp2246 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2247 = (w_sys_tmp2248 + r_run_k_33);
	assign w_sys_tmp2248 = (r_run_copy0_j_65 * w_sys_tmp2245);
	assign w_sys_tmp2250 = (r_run_copy0_j_65 + w_sys_intOne);
	assign w_sys_tmp2251 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp2324 = 32'sh00000020;
	assign w_sys_tmp2325 = ( !w_sys_tmp2326 );
	assign w_sys_tmp2326 = (w_sys_tmp2327 < r_run_j_34);
	assign w_sys_tmp2327 = 32'sh00000031;
	assign w_sys_tmp2329 = (r_run_j_34 - w_sys_tmp2330);
	assign w_sys_tmp2330 = 32'sh0000001f;
	assign w_sys_tmp2332 = (w_sys_tmp2333 + r_run_k_33);
	assign w_sys_tmp2333 = (r_run_tmpj_39 * w_sys_tmp2334);
	assign w_sys_tmp2334 = 32'sh00000081;
	assign w_sys_tmp2335 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2336 = (w_sys_tmp2337 + r_run_k_33);
	assign w_sys_tmp2337 = (r_run_copy0_j_66 * w_sys_tmp2334);
	assign w_sys_tmp2339 = (r_run_copy0_j_66 + w_sys_intOne);
	assign w_sys_tmp2340 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp2413 = 32'sh00000030;
	assign w_sys_tmp2414 = ( !w_sys_tmp2415 );
	assign w_sys_tmp2415 = (w_sys_tmp2416 < r_run_j_34);
	assign w_sys_tmp2416 = 32'sh00000041;
	assign w_sys_tmp2418 = (r_run_j_34 - w_sys_tmp2419);
	assign w_sys_tmp2419 = 32'sh0000002f;
	assign w_sys_tmp2421 = (w_sys_tmp2422 + r_run_k_33);
	assign w_sys_tmp2422 = (r_run_tmpj_39 * w_sys_tmp2423);
	assign w_sys_tmp2423 = 32'sh00000081;
	assign w_sys_tmp2424 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2425 = (w_sys_tmp2426 + r_run_k_33);
	assign w_sys_tmp2426 = (r_run_copy0_j_67 * w_sys_tmp2423);
	assign w_sys_tmp2428 = (r_run_copy0_j_67 + w_sys_intOne);
	assign w_sys_tmp2429 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp2502 = 32'sh00000040;
	assign w_sys_tmp2503 = ( !w_sys_tmp2504 );
	assign w_sys_tmp2504 = (w_sys_tmp2505 < r_run_j_34);
	assign w_sys_tmp2505 = 32'sh00000051;
	assign w_sys_tmp2507 = (r_run_j_34 - w_sys_tmp2508);
	assign w_sys_tmp2508 = 32'sh0000003f;
	assign w_sys_tmp2510 = (w_sys_tmp2511 + r_run_k_33);
	assign w_sys_tmp2511 = (r_run_tmpj_39 * w_sys_tmp2512);
	assign w_sys_tmp2512 = 32'sh00000081;
	assign w_sys_tmp2513 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2514 = (w_sys_tmp2515 + r_run_k_33);
	assign w_sys_tmp2515 = (r_run_copy0_j_68 * w_sys_tmp2512);
	assign w_sys_tmp2517 = (r_run_copy0_j_68 + w_sys_intOne);
	assign w_sys_tmp2518 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp2591 = 32'sh00000050;
	assign w_sys_tmp2592 = ( !w_sys_tmp2593 );
	assign w_sys_tmp2593 = (w_sys_tmp2594 < r_run_j_34);
	assign w_sys_tmp2594 = 32'sh00000061;
	assign w_sys_tmp2596 = (r_run_j_34 - w_sys_tmp2597);
	assign w_sys_tmp2597 = 32'sh0000004f;
	assign w_sys_tmp2599 = (w_sys_tmp2600 + r_run_k_33);
	assign w_sys_tmp2600 = (r_run_tmpj_39 * w_sys_tmp2601);
	assign w_sys_tmp2601 = 32'sh00000081;
	assign w_sys_tmp2602 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2603 = (w_sys_tmp2604 + r_run_k_33);
	assign w_sys_tmp2604 = (r_run_copy0_j_69 * w_sys_tmp2601);
	assign w_sys_tmp2606 = (r_run_copy0_j_69 + w_sys_intOne);
	assign w_sys_tmp2607 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp2680 = 32'sh00000060;
	assign w_sys_tmp2681 = ( !w_sys_tmp2682 );
	assign w_sys_tmp2682 = (w_sys_tmp2683 < r_run_j_34);
	assign w_sys_tmp2683 = 32'sh00000071;
	assign w_sys_tmp2685 = (r_run_j_34 - w_sys_tmp2686);
	assign w_sys_tmp2686 = 32'sh0000005f;
	assign w_sys_tmp2688 = (w_sys_tmp2689 + r_run_k_33);
	assign w_sys_tmp2689 = (r_run_tmpj_39 * w_sys_tmp2690);
	assign w_sys_tmp2690 = 32'sh00000081;
	assign w_sys_tmp2691 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2692 = (w_sys_tmp2693 + r_run_k_33);
	assign w_sys_tmp2693 = (r_run_copy0_j_70 * w_sys_tmp2690);
	assign w_sys_tmp2695 = (r_run_copy0_j_70 + w_sys_intOne);
	assign w_sys_tmp2696 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp2769 = 32'sh00000070;
	assign w_sys_tmp2770 = ( !w_sys_tmp2771 );
	assign w_sys_tmp2771 = (w_sys_tmp2772 < r_run_j_34);
	assign w_sys_tmp2772 = 32'sh00000081;
	assign w_sys_tmp2774 = (r_run_j_34 - w_sys_tmp2775);
	assign w_sys_tmp2775 = 32'sh0000006f;
	assign w_sys_tmp2777 = (w_sys_tmp2778 + r_run_k_33);
	assign w_sys_tmp2778 = (r_run_tmpj_39 * w_sys_tmp2779);
	assign w_sys_tmp2779 = 32'sh00000081;
	assign w_sys_tmp2780 = w_fld_u_0_dataout_1;
	assign w_sys_tmp2781 = (w_sys_tmp2782 + r_run_k_33);
	assign w_sys_tmp2782 = (r_run_copy0_j_71 * w_sys_tmp2779);
	assign w_sys_tmp2784 = (r_run_copy0_j_71 + w_sys_intOne);
	assign w_sys_tmp2785 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp2858 = ( !w_sys_tmp2859 );
	assign w_sys_tmp2859 = (r_run_nlast_38 < r_run_n_35);
	assign w_sys_tmp2860 = (r_run_n_35 + w_sys_intOne);
	assign w_sys_tmp2861 = 32'sh00000002;
	assign w_sys_tmp2862 = ( !w_sys_tmp2863 );
	assign w_sys_tmp2863 = (w_sys_tmp2864 < r_run_k_33);
	assign w_sys_tmp2864 = 32'sh00000020;
	assign w_sys_tmp2867 = (w_sys_tmp2868 + r_run_k_33);
	assign w_sys_tmp2868 = 32'sh00000891;
	assign w_sys_tmp2869 = w_sub01_result_dataout;
	assign w_sys_tmp2870 = (w_sys_tmp2871 + r_run_k_33);
	assign w_sys_tmp2871 = 32'sh00000102;
	assign w_sys_tmp2873 = (w_sys_tmp2874 + r_run_k_33);
	assign w_sys_tmp2874 = 32'sh00000081;
	assign w_sys_tmp2875 = w_sub00_result_dataout;
	assign w_sys_tmp2876 = (w_sys_tmp2877 + r_run_k_33);
	assign w_sys_tmp2877 = 32'sh00000810;
	assign w_sys_tmp2879 = (w_sys_tmp2880 + r_run_k_33);
	assign w_sys_tmp2880 = 32'sh00000912;
	assign w_sys_tmp2897 = w_sub02_result_dataout;
	assign w_sys_tmp2908 = w_sub03_result_dataout;
	assign w_sys_tmp2919 = w_sub04_result_dataout;
	assign w_sys_tmp2930 = w_sub05_result_dataout;
	assign w_sys_tmp2941 = w_sub06_result_dataout;
	assign w_sys_tmp2944 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp2945 = 32'sh00000020;
	assign w_sys_tmp2946 = ( !w_sys_tmp2947 );
	assign w_sys_tmp2947 = (w_sys_tmp2948 < r_run_k_33);
	assign w_sys_tmp2948 = 32'sh00000041;
	assign w_sys_tmp2951 = (w_sys_tmp2952 + r_run_k_33);
	assign w_sys_tmp2952 = 32'sh00000891;
	assign w_sys_tmp2953 = w_sub09_result_dataout;
	assign w_sys_tmp2954 = (w_sys_tmp2955 + r_run_k_33);
	assign w_sys_tmp2955 = 32'sh00000102;
	assign w_sys_tmp2957 = (w_sys_tmp2958 + r_run_k_33);
	assign w_sys_tmp2958 = 32'sh00000081;
	assign w_sys_tmp2959 = w_sub08_result_dataout;
	assign w_sys_tmp2960 = (w_sys_tmp2961 + r_run_k_33);
	assign w_sys_tmp2961 = 32'sh00000810;
	assign w_sys_tmp2963 = (w_sys_tmp2964 + r_run_k_33);
	assign w_sys_tmp2964 = 32'sh00000912;
	assign w_sys_tmp2981 = w_sub10_result_dataout;
	assign w_sys_tmp2992 = w_sub11_result_dataout;
	assign w_sys_tmp3003 = w_sub12_result_dataout;
	assign w_sys_tmp3014 = w_sub13_result_dataout;
	assign w_sys_tmp3025 = w_sub14_result_dataout;
	assign w_sys_tmp3028 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp3029 = 32'sh00000040;
	assign w_sys_tmp3030 = ( !w_sys_tmp3031 );
	assign w_sys_tmp3031 = (w_sys_tmp3032 < r_run_k_33);
	assign w_sys_tmp3032 = 32'sh00000061;
	assign w_sys_tmp3035 = (w_sys_tmp3036 + r_run_k_33);
	assign w_sys_tmp3036 = 32'sh00000891;
	assign w_sys_tmp3037 = w_sub17_result_dataout;
	assign w_sys_tmp3038 = (w_sys_tmp3039 + r_run_k_33);
	assign w_sys_tmp3039 = 32'sh00000102;
	assign w_sys_tmp3041 = (w_sys_tmp3042 + r_run_k_33);
	assign w_sys_tmp3042 = 32'sh00000081;
	assign w_sys_tmp3043 = w_sub16_result_dataout;
	assign w_sys_tmp3044 = (w_sys_tmp3045 + r_run_k_33);
	assign w_sys_tmp3045 = 32'sh00000810;
	assign w_sys_tmp3047 = (w_sys_tmp3048 + r_run_k_33);
	assign w_sys_tmp3048 = 32'sh00000912;
	assign w_sys_tmp3065 = w_sub18_result_dataout;
	assign w_sys_tmp3076 = w_sub19_result_dataout;
	assign w_sys_tmp3087 = w_sub20_result_dataout;
	assign w_sys_tmp3098 = w_sub21_result_dataout;
	assign w_sys_tmp3109 = w_sub22_result_dataout;
	assign w_sys_tmp3112 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp3113 = 32'sh00000060;
	assign w_sys_tmp3114 = ( !w_sys_tmp3115 );
	assign w_sys_tmp3115 = (w_sys_tmp3116 < r_run_k_33);
	assign w_sys_tmp3116 = 32'sh00000081;
	assign w_sys_tmp3119 = (w_sys_tmp3120 + r_run_k_33);
	assign w_sys_tmp3120 = 32'sh00000891;
	assign w_sys_tmp3121 = w_sub25_result_dataout;
	assign w_sys_tmp3122 = (w_sys_tmp3123 + r_run_k_33);
	assign w_sys_tmp3123 = 32'sh00000102;
	assign w_sys_tmp3125 = (w_sys_tmp3126 + r_run_k_33);
	assign w_sys_tmp3126 = 32'sh00000081;
	assign w_sys_tmp3127 = w_sub24_result_dataout;
	assign w_sys_tmp3128 = (w_sys_tmp3129 + r_run_k_33);
	assign w_sys_tmp3129 = 32'sh00000810;
	assign w_sys_tmp3131 = (w_sys_tmp3132 + r_run_k_33);
	assign w_sys_tmp3132 = 32'sh00000912;
	assign w_sys_tmp3149 = w_sub26_result_dataout;
	assign w_sys_tmp3160 = w_sub27_result_dataout;
	assign w_sys_tmp3171 = w_sub28_result_dataout;
	assign w_sys_tmp3182 = w_sub29_result_dataout;
	assign w_sys_tmp3193 = w_sub30_result_dataout;
	assign w_sys_tmp3196 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp3197 = ( !w_sys_tmp3198 );
	assign w_sys_tmp3198 = (w_sys_tmp3199 < r_run_j_34);
	assign w_sys_tmp3199 = 32'sh00000011;
	assign w_sys_tmp3202 = (w_sys_tmp3203 + w_sys_tmp3205);
	assign w_sys_tmp3203 = (r_run_j_34 * w_sys_tmp3204);
	assign w_sys_tmp3204 = 32'sh00000081;
	assign w_sys_tmp3205 = 32'sh00000021;
	assign w_sys_tmp3206 = w_sub08_result_dataout;
	assign w_sys_tmp3207 = (w_sys_tmp3208 + w_sys_tmp3205);
	assign w_sys_tmp3208 = (r_run_copy10_j_82 * w_sys_tmp3204);
	assign w_sys_tmp3212 = (w_sys_tmp3213 + w_sys_tmp3215);
	assign w_sys_tmp3213 = (r_run_copy9_j_81 * w_sys_tmp3204);
	assign w_sys_tmp3215 = 32'sh00000020;
	assign w_sys_tmp3216 = w_sub00_result_dataout;
	assign w_sys_tmp3217 = (w_sys_tmp3218 + w_sys_tmp3215);
	assign w_sys_tmp3218 = (r_run_copy8_j_80 * w_sys_tmp3204);
	assign w_sys_tmp3222 = (w_sys_tmp3223 + w_sys_tmp3225);
	assign w_sys_tmp3223 = (r_run_copy7_j_79 * w_sys_tmp3204);
	assign w_sys_tmp3225 = 32'sh00000041;
	assign w_sys_tmp3226 = (w_sys_tmp3227 + w_sys_tmp3225);
	assign w_sys_tmp3227 = (r_run_copy6_j_78 * w_sys_tmp3204);
	assign w_sys_tmp3231 = (w_sys_tmp3232 + w_sys_tmp3234);
	assign w_sys_tmp3232 = (r_run_copy5_j_77 * w_sys_tmp3204);
	assign w_sys_tmp3234 = 32'sh00000040;
	assign w_sys_tmp3236 = (w_sys_tmp3237 + w_sys_tmp3234);
	assign w_sys_tmp3237 = (r_run_copy4_j_76 * w_sys_tmp3204);
	assign w_sys_tmp3241 = (w_sys_tmp3242 + w_sys_tmp3244);
	assign w_sys_tmp3242 = (r_run_copy3_j_75 * w_sys_tmp3204);
	assign w_sys_tmp3244 = 32'sh00000061;
	assign w_sys_tmp3245 = (w_sys_tmp3246 + w_sys_tmp3244);
	assign w_sys_tmp3246 = (r_run_copy2_j_74 * w_sys_tmp3204);
	assign w_sys_tmp3250 = (w_sys_tmp3251 + w_sys_tmp3253);
	assign w_sys_tmp3251 = (r_run_copy1_j_73 * w_sys_tmp3204);
	assign w_sys_tmp3253 = 32'sh00000060;
	assign w_sys_tmp3254 = w_sub16_result_dataout;
	assign w_sys_tmp3255 = (w_sys_tmp3256 + w_sys_tmp3253);
	assign w_sys_tmp3256 = (r_run_copy0_j_72 * w_sys_tmp3204);
	assign w_sys_tmp3259 = (r_run_copy0_j_72 + w_sys_intOne);
	assign w_sys_tmp3260 = (r_run_copy1_j_73 + w_sys_intOne);
	assign w_sys_tmp3261 = (r_run_copy2_j_74 + w_sys_intOne);
	assign w_sys_tmp3262 = (r_run_copy3_j_75 + w_sys_intOne);
	assign w_sys_tmp3263 = (r_run_copy4_j_76 + w_sys_intOne);
	assign w_sys_tmp3264 = (r_run_copy5_j_77 + w_sys_intOne);
	assign w_sys_tmp3265 = (r_run_copy6_j_78 + w_sys_intOne);
	assign w_sys_tmp3266 = (r_run_copy7_j_79 + w_sys_intOne);
	assign w_sys_tmp3267 = (r_run_copy8_j_80 + w_sys_intOne);
	assign w_sys_tmp3268 = (r_run_copy9_j_81 + w_sys_intOne);
	assign w_sys_tmp3269 = (r_run_copy10_j_82 + w_sys_intOne);
	assign w_sys_tmp3270 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp3697 = 32'sh00000010;
	assign w_sys_tmp3698 = ( !w_sys_tmp3699 );
	assign w_sys_tmp3699 = (w_sys_tmp3700 < r_run_j_34);
	assign w_sys_tmp3700 = 32'sh00000021;
	assign w_sys_tmp3703 = (w_sys_tmp3704 + w_sys_tmp3706);
	assign w_sys_tmp3704 = (r_run_j_34 * w_sys_tmp3705);
	assign w_sys_tmp3705 = 32'sh00000081;
	assign w_sys_tmp3706 = 32'sh00000021;
	assign w_sys_tmp3707 = w_sub09_result_dataout;
	assign w_sys_tmp3708 = (w_sys_tmp3709 + w_sys_tmp3706);
	assign w_sys_tmp3709 = (r_run_copy10_j_93 * w_sys_tmp3705);
	assign w_sys_tmp3713 = (w_sys_tmp3714 + w_sys_tmp3716);
	assign w_sys_tmp3714 = (r_run_copy9_j_92 * w_sys_tmp3705);
	assign w_sys_tmp3716 = 32'sh00000020;
	assign w_sys_tmp3717 = w_sub01_result_dataout;
	assign w_sys_tmp3718 = (w_sys_tmp3719 + w_sys_tmp3716);
	assign w_sys_tmp3719 = (r_run_copy8_j_91 * w_sys_tmp3705);
	assign w_sys_tmp3723 = (w_sys_tmp3724 + w_sys_tmp3726);
	assign w_sys_tmp3724 = (r_run_copy7_j_90 * w_sys_tmp3705);
	assign w_sys_tmp3726 = 32'sh00000041;
	assign w_sys_tmp3727 = (w_sys_tmp3728 + w_sys_tmp3726);
	assign w_sys_tmp3728 = (r_run_copy6_j_89 * w_sys_tmp3705);
	assign w_sys_tmp3732 = (w_sys_tmp3733 + w_sys_tmp3735);
	assign w_sys_tmp3733 = (r_run_copy5_j_88 * w_sys_tmp3705);
	assign w_sys_tmp3735 = 32'sh00000040;
	assign w_sys_tmp3737 = (w_sys_tmp3738 + w_sys_tmp3735);
	assign w_sys_tmp3738 = (r_run_copy4_j_87 * w_sys_tmp3705);
	assign w_sys_tmp3742 = (w_sys_tmp3743 + w_sys_tmp3745);
	assign w_sys_tmp3743 = (r_run_copy3_j_86 * w_sys_tmp3705);
	assign w_sys_tmp3745 = 32'sh00000061;
	assign w_sys_tmp3746 = (w_sys_tmp3747 + w_sys_tmp3745);
	assign w_sys_tmp3747 = (r_run_copy2_j_85 * w_sys_tmp3705);
	assign w_sys_tmp3751 = (w_sys_tmp3752 + w_sys_tmp3754);
	assign w_sys_tmp3752 = (r_run_copy1_j_84 * w_sys_tmp3705);
	assign w_sys_tmp3754 = 32'sh00000060;
	assign w_sys_tmp3755 = w_sub17_result_dataout;
	assign w_sys_tmp3756 = (w_sys_tmp3757 + w_sys_tmp3754);
	assign w_sys_tmp3757 = (r_run_copy0_j_83 * w_sys_tmp3705);
	assign w_sys_tmp3760 = (r_run_copy0_j_83 + w_sys_intOne);
	assign w_sys_tmp3761 = (r_run_copy1_j_84 + w_sys_intOne);
	assign w_sys_tmp3762 = (r_run_copy2_j_85 + w_sys_intOne);
	assign w_sys_tmp3763 = (r_run_copy3_j_86 + w_sys_intOne);
	assign w_sys_tmp3764 = (r_run_copy4_j_87 + w_sys_intOne);
	assign w_sys_tmp3765 = (r_run_copy5_j_88 + w_sys_intOne);
	assign w_sys_tmp3766 = (r_run_copy6_j_89 + w_sys_intOne);
	assign w_sys_tmp3767 = (r_run_copy7_j_90 + w_sys_intOne);
	assign w_sys_tmp3768 = (r_run_copy8_j_91 + w_sys_intOne);
	assign w_sys_tmp3769 = (r_run_copy9_j_92 + w_sys_intOne);
	assign w_sys_tmp3770 = (r_run_copy10_j_93 + w_sys_intOne);
	assign w_sys_tmp3771 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp4198 = 32'sh00000020;
	assign w_sys_tmp4199 = ( !w_sys_tmp4200 );
	assign w_sys_tmp4200 = (w_sys_tmp4201 < r_run_j_34);
	assign w_sys_tmp4201 = 32'sh00000031;
	assign w_sys_tmp4204 = (w_sys_tmp4205 + w_sys_tmp4207);
	assign w_sys_tmp4205 = (r_run_j_34 * w_sys_tmp4206);
	assign w_sys_tmp4206 = 32'sh00000081;
	assign w_sys_tmp4207 = 32'sh00000021;
	assign w_sys_tmp4208 = w_sub10_result_dataout;
	assign w_sys_tmp4209 = (w_sys_tmp4210 + w_sys_tmp4207);
	assign w_sys_tmp4210 = (r_run_copy10_j_104 * w_sys_tmp4206);
	assign w_sys_tmp4214 = (w_sys_tmp4215 + w_sys_tmp4217);
	assign w_sys_tmp4215 = (r_run_copy9_j_103 * w_sys_tmp4206);
	assign w_sys_tmp4217 = 32'sh00000020;
	assign w_sys_tmp4218 = w_sub02_result_dataout;
	assign w_sys_tmp4219 = (w_sys_tmp4220 + w_sys_tmp4217);
	assign w_sys_tmp4220 = (r_run_copy8_j_102 * w_sys_tmp4206);
	assign w_sys_tmp4224 = (w_sys_tmp4225 + w_sys_tmp4227);
	assign w_sys_tmp4225 = (r_run_copy7_j_101 * w_sys_tmp4206);
	assign w_sys_tmp4227 = 32'sh00000041;
	assign w_sys_tmp4228 = (w_sys_tmp4229 + w_sys_tmp4227);
	assign w_sys_tmp4229 = (r_run_copy6_j_100 * w_sys_tmp4206);
	assign w_sys_tmp4233 = (w_sys_tmp4234 + w_sys_tmp4236);
	assign w_sys_tmp4234 = (r_run_copy5_j_99 * w_sys_tmp4206);
	assign w_sys_tmp4236 = 32'sh00000040;
	assign w_sys_tmp4238 = (w_sys_tmp4239 + w_sys_tmp4236);
	assign w_sys_tmp4239 = (r_run_copy4_j_98 * w_sys_tmp4206);
	assign w_sys_tmp4243 = (w_sys_tmp4244 + w_sys_tmp4246);
	assign w_sys_tmp4244 = (r_run_copy3_j_97 * w_sys_tmp4206);
	assign w_sys_tmp4246 = 32'sh00000061;
	assign w_sys_tmp4247 = (w_sys_tmp4248 + w_sys_tmp4246);
	assign w_sys_tmp4248 = (r_run_copy2_j_96 * w_sys_tmp4206);
	assign w_sys_tmp4252 = (w_sys_tmp4253 + w_sys_tmp4255);
	assign w_sys_tmp4253 = (r_run_copy1_j_95 * w_sys_tmp4206);
	assign w_sys_tmp4255 = 32'sh00000060;
	assign w_sys_tmp4256 = w_sub18_result_dataout;
	assign w_sys_tmp4257 = (w_sys_tmp4258 + w_sys_tmp4255);
	assign w_sys_tmp4258 = (r_run_copy0_j_94 * w_sys_tmp4206);
	assign w_sys_tmp4261 = (r_run_copy0_j_94 + w_sys_intOne);
	assign w_sys_tmp4262 = (r_run_copy1_j_95 + w_sys_intOne);
	assign w_sys_tmp4263 = (r_run_copy2_j_96 + w_sys_intOne);
	assign w_sys_tmp4264 = (r_run_copy3_j_97 + w_sys_intOne);
	assign w_sys_tmp4265 = (r_run_copy4_j_98 + w_sys_intOne);
	assign w_sys_tmp4266 = (r_run_copy5_j_99 + w_sys_intOne);
	assign w_sys_tmp4267 = (r_run_copy6_j_100 + w_sys_intOne);
	assign w_sys_tmp4268 = (r_run_copy7_j_101 + w_sys_intOne);
	assign w_sys_tmp4269 = (r_run_copy8_j_102 + w_sys_intOne);
	assign w_sys_tmp4270 = (r_run_copy9_j_103 + w_sys_intOne);
	assign w_sys_tmp4271 = (r_run_copy10_j_104 + w_sys_intOne);
	assign w_sys_tmp4272 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp4699 = 32'sh00000030;
	assign w_sys_tmp4700 = ( !w_sys_tmp4701 );
	assign w_sys_tmp4701 = (w_sys_tmp4702 < r_run_j_34);
	assign w_sys_tmp4702 = 32'sh00000041;
	assign w_sys_tmp4705 = (w_sys_tmp4706 + w_sys_tmp4708);
	assign w_sys_tmp4706 = (r_run_j_34 * w_sys_tmp4707);
	assign w_sys_tmp4707 = 32'sh00000081;
	assign w_sys_tmp4708 = 32'sh00000021;
	assign w_sys_tmp4709 = w_sub11_result_dataout;
	assign w_sys_tmp4710 = (w_sys_tmp4711 + w_sys_tmp4708);
	assign w_sys_tmp4711 = (r_run_copy10_j_115 * w_sys_tmp4707);
	assign w_sys_tmp4715 = (w_sys_tmp4716 + w_sys_tmp4718);
	assign w_sys_tmp4716 = (r_run_copy9_j_114 * w_sys_tmp4707);
	assign w_sys_tmp4718 = 32'sh00000020;
	assign w_sys_tmp4719 = w_sub03_result_dataout;
	assign w_sys_tmp4720 = (w_sys_tmp4721 + w_sys_tmp4718);
	assign w_sys_tmp4721 = (r_run_copy8_j_113 * w_sys_tmp4707);
	assign w_sys_tmp4725 = (w_sys_tmp4726 + w_sys_tmp4728);
	assign w_sys_tmp4726 = (r_run_copy7_j_112 * w_sys_tmp4707);
	assign w_sys_tmp4728 = 32'sh00000041;
	assign w_sys_tmp4729 = (w_sys_tmp4730 + w_sys_tmp4728);
	assign w_sys_tmp4730 = (r_run_copy6_j_111 * w_sys_tmp4707);
	assign w_sys_tmp4734 = (w_sys_tmp4735 + w_sys_tmp4737);
	assign w_sys_tmp4735 = (r_run_copy5_j_110 * w_sys_tmp4707);
	assign w_sys_tmp4737 = 32'sh00000040;
	assign w_sys_tmp4739 = (w_sys_tmp4740 + w_sys_tmp4737);
	assign w_sys_tmp4740 = (r_run_copy4_j_109 * w_sys_tmp4707);
	assign w_sys_tmp4744 = (w_sys_tmp4745 + w_sys_tmp4747);
	assign w_sys_tmp4745 = (r_run_copy3_j_108 * w_sys_tmp4707);
	assign w_sys_tmp4747 = 32'sh00000061;
	assign w_sys_tmp4748 = (w_sys_tmp4749 + w_sys_tmp4747);
	assign w_sys_tmp4749 = (r_run_copy2_j_107 * w_sys_tmp4707);
	assign w_sys_tmp4753 = (w_sys_tmp4754 + w_sys_tmp4756);
	assign w_sys_tmp4754 = (r_run_copy1_j_106 * w_sys_tmp4707);
	assign w_sys_tmp4756 = 32'sh00000060;
	assign w_sys_tmp4757 = w_sub19_result_dataout;
	assign w_sys_tmp4758 = (w_sys_tmp4759 + w_sys_tmp4756);
	assign w_sys_tmp4759 = (r_run_copy0_j_105 * w_sys_tmp4707);
	assign w_sys_tmp4762 = (r_run_copy0_j_105 + w_sys_intOne);
	assign w_sys_tmp4763 = (r_run_copy1_j_106 + w_sys_intOne);
	assign w_sys_tmp4764 = (r_run_copy2_j_107 + w_sys_intOne);
	assign w_sys_tmp4765 = (r_run_copy3_j_108 + w_sys_intOne);
	assign w_sys_tmp4766 = (r_run_copy4_j_109 + w_sys_intOne);
	assign w_sys_tmp4767 = (r_run_copy5_j_110 + w_sys_intOne);
	assign w_sys_tmp4768 = (r_run_copy6_j_111 + w_sys_intOne);
	assign w_sys_tmp4769 = (r_run_copy7_j_112 + w_sys_intOne);
	assign w_sys_tmp4770 = (r_run_copy8_j_113 + w_sys_intOne);
	assign w_sys_tmp4771 = (r_run_copy9_j_114 + w_sys_intOne);
	assign w_sys_tmp4772 = (r_run_copy10_j_115 + w_sys_intOne);
	assign w_sys_tmp4773 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp5200 = 32'sh00000040;
	assign w_sys_tmp5201 = ( !w_sys_tmp5202 );
	assign w_sys_tmp5202 = (w_sys_tmp5203 < r_run_j_34);
	assign w_sys_tmp5203 = 32'sh00000051;
	assign w_sys_tmp5206 = (w_sys_tmp5207 + w_sys_tmp5209);
	assign w_sys_tmp5207 = (r_run_j_34 * w_sys_tmp5208);
	assign w_sys_tmp5208 = 32'sh00000081;
	assign w_sys_tmp5209 = 32'sh00000021;
	assign w_sys_tmp5210 = w_sub12_result_dataout;
	assign w_sys_tmp5211 = (w_sys_tmp5212 + w_sys_tmp5209);
	assign w_sys_tmp5212 = (r_run_copy10_j_126 * w_sys_tmp5208);
	assign w_sys_tmp5216 = (w_sys_tmp5217 + w_sys_tmp5219);
	assign w_sys_tmp5217 = (r_run_copy9_j_125 * w_sys_tmp5208);
	assign w_sys_tmp5219 = 32'sh00000020;
	assign w_sys_tmp5220 = w_sub04_result_dataout;
	assign w_sys_tmp5221 = (w_sys_tmp5222 + w_sys_tmp5219);
	assign w_sys_tmp5222 = (r_run_copy8_j_124 * w_sys_tmp5208);
	assign w_sys_tmp5226 = (w_sys_tmp5227 + w_sys_tmp5229);
	assign w_sys_tmp5227 = (r_run_copy7_j_123 * w_sys_tmp5208);
	assign w_sys_tmp5229 = 32'sh00000041;
	assign w_sys_tmp5230 = (w_sys_tmp5231 + w_sys_tmp5229);
	assign w_sys_tmp5231 = (r_run_copy6_j_122 * w_sys_tmp5208);
	assign w_sys_tmp5235 = (w_sys_tmp5236 + w_sys_tmp5238);
	assign w_sys_tmp5236 = (r_run_copy5_j_121 * w_sys_tmp5208);
	assign w_sys_tmp5238 = 32'sh00000040;
	assign w_sys_tmp5240 = (w_sys_tmp5241 + w_sys_tmp5238);
	assign w_sys_tmp5241 = (r_run_copy4_j_120 * w_sys_tmp5208);
	assign w_sys_tmp5245 = (w_sys_tmp5246 + w_sys_tmp5248);
	assign w_sys_tmp5246 = (r_run_copy3_j_119 * w_sys_tmp5208);
	assign w_sys_tmp5248 = 32'sh00000061;
	assign w_sys_tmp5249 = (w_sys_tmp5250 + w_sys_tmp5248);
	assign w_sys_tmp5250 = (r_run_copy2_j_118 * w_sys_tmp5208);
	assign w_sys_tmp5254 = (w_sys_tmp5255 + w_sys_tmp5257);
	assign w_sys_tmp5255 = (r_run_copy1_j_117 * w_sys_tmp5208);
	assign w_sys_tmp5257 = 32'sh00000060;
	assign w_sys_tmp5258 = w_sub20_result_dataout;
	assign w_sys_tmp5259 = (w_sys_tmp5260 + w_sys_tmp5257);
	assign w_sys_tmp5260 = (r_run_copy0_j_116 * w_sys_tmp5208);
	assign w_sys_tmp5263 = (r_run_copy0_j_116 + w_sys_intOne);
	assign w_sys_tmp5264 = (r_run_copy1_j_117 + w_sys_intOne);
	assign w_sys_tmp5265 = (r_run_copy2_j_118 + w_sys_intOne);
	assign w_sys_tmp5266 = (r_run_copy3_j_119 + w_sys_intOne);
	assign w_sys_tmp5267 = (r_run_copy4_j_120 + w_sys_intOne);
	assign w_sys_tmp5268 = (r_run_copy5_j_121 + w_sys_intOne);
	assign w_sys_tmp5269 = (r_run_copy6_j_122 + w_sys_intOne);
	assign w_sys_tmp5270 = (r_run_copy7_j_123 + w_sys_intOne);
	assign w_sys_tmp5271 = (r_run_copy8_j_124 + w_sys_intOne);
	assign w_sys_tmp5272 = (r_run_copy9_j_125 + w_sys_intOne);
	assign w_sys_tmp5273 = (r_run_copy10_j_126 + w_sys_intOne);
	assign w_sys_tmp5274 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp5701 = 32'sh00000050;
	assign w_sys_tmp5702 = ( !w_sys_tmp5703 );
	assign w_sys_tmp5703 = (w_sys_tmp5704 < r_run_j_34);
	assign w_sys_tmp5704 = 32'sh00000061;
	assign w_sys_tmp5707 = (w_sys_tmp5708 + w_sys_tmp5710);
	assign w_sys_tmp5708 = (r_run_j_34 * w_sys_tmp5709);
	assign w_sys_tmp5709 = 32'sh00000081;
	assign w_sys_tmp5710 = 32'sh00000021;
	assign w_sys_tmp5711 = w_sub13_result_dataout;
	assign w_sys_tmp5712 = (w_sys_tmp5713 + w_sys_tmp5710);
	assign w_sys_tmp5713 = (r_run_copy10_j_137 * w_sys_tmp5709);
	assign w_sys_tmp5717 = (w_sys_tmp5718 + w_sys_tmp5720);
	assign w_sys_tmp5718 = (r_run_copy9_j_136 * w_sys_tmp5709);
	assign w_sys_tmp5720 = 32'sh00000020;
	assign w_sys_tmp5721 = w_sub05_result_dataout;
	assign w_sys_tmp5722 = (w_sys_tmp5723 + w_sys_tmp5720);
	assign w_sys_tmp5723 = (r_run_copy8_j_135 * w_sys_tmp5709);
	assign w_sys_tmp5727 = (w_sys_tmp5728 + w_sys_tmp5730);
	assign w_sys_tmp5728 = (r_run_copy7_j_134 * w_sys_tmp5709);
	assign w_sys_tmp5730 = 32'sh00000041;
	assign w_sys_tmp5731 = (w_sys_tmp5732 + w_sys_tmp5730);
	assign w_sys_tmp5732 = (r_run_copy6_j_133 * w_sys_tmp5709);
	assign w_sys_tmp5736 = (w_sys_tmp5737 + w_sys_tmp5739);
	assign w_sys_tmp5737 = (r_run_copy5_j_132 * w_sys_tmp5709);
	assign w_sys_tmp5739 = 32'sh00000040;
	assign w_sys_tmp5741 = (w_sys_tmp5742 + w_sys_tmp5739);
	assign w_sys_tmp5742 = (r_run_copy4_j_131 * w_sys_tmp5709);
	assign w_sys_tmp5746 = (w_sys_tmp5747 + w_sys_tmp5749);
	assign w_sys_tmp5747 = (r_run_copy3_j_130 * w_sys_tmp5709);
	assign w_sys_tmp5749 = 32'sh00000061;
	assign w_sys_tmp5750 = (w_sys_tmp5751 + w_sys_tmp5749);
	assign w_sys_tmp5751 = (r_run_copy2_j_129 * w_sys_tmp5709);
	assign w_sys_tmp5755 = (w_sys_tmp5756 + w_sys_tmp5758);
	assign w_sys_tmp5756 = (r_run_copy1_j_128 * w_sys_tmp5709);
	assign w_sys_tmp5758 = 32'sh00000060;
	assign w_sys_tmp5759 = w_sub21_result_dataout;
	assign w_sys_tmp5760 = (w_sys_tmp5761 + w_sys_tmp5758);
	assign w_sys_tmp5761 = (r_run_copy0_j_127 * w_sys_tmp5709);
	assign w_sys_tmp5764 = (r_run_copy0_j_127 + w_sys_intOne);
	assign w_sys_tmp5765 = (r_run_copy1_j_128 + w_sys_intOne);
	assign w_sys_tmp5766 = (r_run_copy2_j_129 + w_sys_intOne);
	assign w_sys_tmp5767 = (r_run_copy3_j_130 + w_sys_intOne);
	assign w_sys_tmp5768 = (r_run_copy4_j_131 + w_sys_intOne);
	assign w_sys_tmp5769 = (r_run_copy5_j_132 + w_sys_intOne);
	assign w_sys_tmp5770 = (r_run_copy6_j_133 + w_sys_intOne);
	assign w_sys_tmp5771 = (r_run_copy7_j_134 + w_sys_intOne);
	assign w_sys_tmp5772 = (r_run_copy8_j_135 + w_sys_intOne);
	assign w_sys_tmp5773 = (r_run_copy9_j_136 + w_sys_intOne);
	assign w_sys_tmp5774 = (r_run_copy10_j_137 + w_sys_intOne);
	assign w_sys_tmp5775 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp6202 = 32'sh00000060;
	assign w_sys_tmp6203 = ( !w_sys_tmp6204 );
	assign w_sys_tmp6204 = (w_sys_tmp6205 < r_run_j_34);
	assign w_sys_tmp6205 = 32'sh00000071;
	assign w_sys_tmp6208 = (w_sys_tmp6209 + w_sys_tmp6211);
	assign w_sys_tmp6209 = (r_run_j_34 * w_sys_tmp6210);
	assign w_sys_tmp6210 = 32'sh00000081;
	assign w_sys_tmp6211 = 32'sh00000021;
	assign w_sys_tmp6212 = w_sub14_result_dataout;
	assign w_sys_tmp6213 = (w_sys_tmp6214 + w_sys_tmp6211);
	assign w_sys_tmp6214 = (r_run_copy10_j_148 * w_sys_tmp6210);
	assign w_sys_tmp6218 = (w_sys_tmp6219 + w_sys_tmp6221);
	assign w_sys_tmp6219 = (r_run_copy9_j_147 * w_sys_tmp6210);
	assign w_sys_tmp6221 = 32'sh00000020;
	assign w_sys_tmp6222 = w_sub06_result_dataout;
	assign w_sys_tmp6223 = (w_sys_tmp6224 + w_sys_tmp6221);
	assign w_sys_tmp6224 = (r_run_copy8_j_146 * w_sys_tmp6210);
	assign w_sys_tmp6228 = (w_sys_tmp6229 + w_sys_tmp6231);
	assign w_sys_tmp6229 = (r_run_copy7_j_145 * w_sys_tmp6210);
	assign w_sys_tmp6231 = 32'sh00000041;
	assign w_sys_tmp6232 = (w_sys_tmp6233 + w_sys_tmp6231);
	assign w_sys_tmp6233 = (r_run_copy6_j_144 * w_sys_tmp6210);
	assign w_sys_tmp6237 = (w_sys_tmp6238 + w_sys_tmp6240);
	assign w_sys_tmp6238 = (r_run_copy5_j_143 * w_sys_tmp6210);
	assign w_sys_tmp6240 = 32'sh00000040;
	assign w_sys_tmp6242 = (w_sys_tmp6243 + w_sys_tmp6240);
	assign w_sys_tmp6243 = (r_run_copy4_j_142 * w_sys_tmp6210);
	assign w_sys_tmp6247 = (w_sys_tmp6248 + w_sys_tmp6250);
	assign w_sys_tmp6248 = (r_run_copy3_j_141 * w_sys_tmp6210);
	assign w_sys_tmp6250 = 32'sh00000061;
	assign w_sys_tmp6251 = (w_sys_tmp6252 + w_sys_tmp6250);
	assign w_sys_tmp6252 = (r_run_copy2_j_140 * w_sys_tmp6210);
	assign w_sys_tmp6256 = (w_sys_tmp6257 + w_sys_tmp6259);
	assign w_sys_tmp6257 = (r_run_copy1_j_139 * w_sys_tmp6210);
	assign w_sys_tmp6259 = 32'sh00000060;
	assign w_sys_tmp6260 = w_sub22_result_dataout;
	assign w_sys_tmp6261 = (w_sys_tmp6262 + w_sys_tmp6259);
	assign w_sys_tmp6262 = (r_run_copy0_j_138 * w_sys_tmp6210);
	assign w_sys_tmp6265 = (r_run_copy0_j_138 + w_sys_intOne);
	assign w_sys_tmp6266 = (r_run_copy1_j_139 + w_sys_intOne);
	assign w_sys_tmp6267 = (r_run_copy2_j_140 + w_sys_intOne);
	assign w_sys_tmp6268 = (r_run_copy3_j_141 + w_sys_intOne);
	assign w_sys_tmp6269 = (r_run_copy4_j_142 + w_sys_intOne);
	assign w_sys_tmp6270 = (r_run_copy5_j_143 + w_sys_intOne);
	assign w_sys_tmp6271 = (r_run_copy6_j_144 + w_sys_intOne);
	assign w_sys_tmp6272 = (r_run_copy7_j_145 + w_sys_intOne);
	assign w_sys_tmp6273 = (r_run_copy8_j_146 + w_sys_intOne);
	assign w_sys_tmp6274 = (r_run_copy9_j_147 + w_sys_intOne);
	assign w_sys_tmp6275 = (r_run_copy10_j_148 + w_sys_intOne);
	assign w_sys_tmp6276 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp6703 = 32'sh00000070;
	assign w_sys_tmp6704 = ( !w_sys_tmp6705 );
	assign w_sys_tmp6705 = (w_sys_tmp6706 < r_run_j_34);
	assign w_sys_tmp6706 = 32'sh00000081;
	assign w_sys_tmp6709 = (w_sys_tmp6710 + w_sys_tmp6712);
	assign w_sys_tmp6710 = (r_run_j_34 * w_sys_tmp6711);
	assign w_sys_tmp6711 = 32'sh00000081;
	assign w_sys_tmp6712 = 32'sh00000021;
	assign w_sys_tmp6713 = w_sub15_result_dataout;
	assign w_sys_tmp6714 = (w_sys_tmp6715 + w_sys_tmp6712);
	assign w_sys_tmp6715 = (r_run_copy10_j_159 * w_sys_tmp6711);
	assign w_sys_tmp6719 = (w_sys_tmp6720 + w_sys_tmp6722);
	assign w_sys_tmp6720 = (r_run_copy9_j_158 * w_sys_tmp6711);
	assign w_sys_tmp6722 = 32'sh00000020;
	assign w_sys_tmp6723 = w_sub07_result_dataout;
	assign w_sys_tmp6724 = (w_sys_tmp6725 + w_sys_tmp6722);
	assign w_sys_tmp6725 = (r_run_copy8_j_157 * w_sys_tmp6711);
	assign w_sys_tmp6729 = (w_sys_tmp6730 + w_sys_tmp6732);
	assign w_sys_tmp6730 = (r_run_copy7_j_156 * w_sys_tmp6711);
	assign w_sys_tmp6732 = 32'sh00000041;
	assign w_sys_tmp6733 = (w_sys_tmp6734 + w_sys_tmp6732);
	assign w_sys_tmp6734 = (r_run_copy6_j_155 * w_sys_tmp6711);
	assign w_sys_tmp6738 = (w_sys_tmp6739 + w_sys_tmp6741);
	assign w_sys_tmp6739 = (r_run_copy5_j_154 * w_sys_tmp6711);
	assign w_sys_tmp6741 = 32'sh00000040;
	assign w_sys_tmp6743 = (w_sys_tmp6744 + w_sys_tmp6741);
	assign w_sys_tmp6744 = (r_run_copy4_j_153 * w_sys_tmp6711);
	assign w_sys_tmp6748 = (w_sys_tmp6749 + w_sys_tmp6751);
	assign w_sys_tmp6749 = (r_run_copy3_j_152 * w_sys_tmp6711);
	assign w_sys_tmp6751 = 32'sh00000061;
	assign w_sys_tmp6752 = (w_sys_tmp6753 + w_sys_tmp6751);
	assign w_sys_tmp6753 = (r_run_copy2_j_151 * w_sys_tmp6711);
	assign w_sys_tmp6757 = (w_sys_tmp6758 + w_sys_tmp6760);
	assign w_sys_tmp6758 = (r_run_copy1_j_150 * w_sys_tmp6711);
	assign w_sys_tmp6760 = 32'sh00000060;
	assign w_sys_tmp6761 = w_sub16_result_dataout;
	assign w_sys_tmp6762 = (w_sys_tmp6763 + w_sys_tmp6760);
	assign w_sys_tmp6763 = (r_run_copy0_j_149 * w_sys_tmp6711);
	assign w_sys_tmp6766 = (r_run_copy0_j_149 + w_sys_intOne);
	assign w_sys_tmp6767 = (r_run_copy1_j_150 + w_sys_intOne);
	assign w_sys_tmp6768 = (r_run_copy2_j_151 + w_sys_intOne);
	assign w_sys_tmp6769 = (r_run_copy3_j_152 + w_sys_intOne);
	assign w_sys_tmp6770 = (r_run_copy4_j_153 + w_sys_intOne);
	assign w_sys_tmp6771 = (r_run_copy5_j_154 + w_sys_intOne);
	assign w_sys_tmp6772 = (r_run_copy6_j_155 + w_sys_intOne);
	assign w_sys_tmp6773 = (r_run_copy7_j_156 + w_sys_intOne);
	assign w_sys_tmp6774 = (r_run_copy8_j_157 + w_sys_intOne);
	assign w_sys_tmp6775 = (r_run_copy9_j_158 + w_sys_intOne);
	assign w_sys_tmp6776 = (r_run_copy10_j_159 + w_sys_intOne);
	assign w_sys_tmp6777 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp7192 = 32'sh00000002;
	assign w_sys_tmp7193 = ( !w_sys_tmp7194 );
	assign w_sys_tmp7194 = (w_sys_tmp7195 < r_run_k_33);
	assign w_sys_tmp7195 = 32'sh00000020;
	assign w_sys_tmp7196 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp7197 = 32'sh00000002;
	assign w_sys_tmp7198 = ( !w_sys_tmp7199 );
	assign w_sys_tmp7199 = (w_sys_tmp7200 < r_run_j_34);
	assign w_sys_tmp7200 = 32'sh00000010;
	assign w_sys_tmp7203 = (w_sys_tmp7204 + r_run_k_33);
	assign w_sys_tmp7204 = (r_run_j_34 * w_sys_tmp7205);
	assign w_sys_tmp7205 = 32'sh00000081;
	assign w_sys_tmp7206 = w_sub00_result_dataout;
	assign w_sys_tmp7207 = (w_sys_tmp7208 + r_run_k_33);
	assign w_sys_tmp7208 = (r_run_copy0_j_160 * w_sys_tmp7205);
	assign w_sys_tmp7210 = (r_run_copy0_j_160 + w_sys_intOne);
	assign w_sys_tmp7211 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp7272 = 32'sh00000011;
	assign w_sys_tmp7273 = ( !w_sys_tmp7274 );
	assign w_sys_tmp7274 = (w_sys_tmp7275 < r_run_j_34);
	assign w_sys_tmp7275 = 32'sh00000020;
	assign w_sys_tmp7277 = (r_run_j_34 - w_sys_tmp7278);
	assign w_sys_tmp7278 = 32'sh0000000f;
	assign w_sys_tmp7280 = (w_sys_tmp7281 + r_run_k_33);
	assign w_sys_tmp7281 = (r_run_copy1_j_162 * w_sys_tmp7282);
	assign w_sys_tmp7282 = 32'sh00000081;
	assign w_sys_tmp7283 = w_sub01_result_dataout;
	assign w_sys_tmp7284 = (w_sys_tmp7285 + r_run_k_33);
	assign w_sys_tmp7285 = (r_run_copy0_j_161 * w_sys_tmp7282);
	assign w_sys_tmp7287 = (r_run_copy0_j_161 + w_sys_intOne);
	assign w_sys_tmp7288 = (r_run_copy1_j_162 + w_sys_intOne);
	assign w_sys_tmp7289 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp7368 = 32'sh00000021;
	assign w_sys_tmp7369 = ( !w_sys_tmp7370 );
	assign w_sys_tmp7370 = (w_sys_tmp7371 < r_run_j_34);
	assign w_sys_tmp7371 = 32'sh00000030;
	assign w_sys_tmp7373 = (r_run_j_34 - w_sys_tmp7374);
	assign w_sys_tmp7374 = 32'sh0000001f;
	assign w_sys_tmp7376 = (w_sys_tmp7377 + r_run_k_33);
	assign w_sys_tmp7377 = (r_run_copy1_j_164 * w_sys_tmp7378);
	assign w_sys_tmp7378 = 32'sh00000081;
	assign w_sys_tmp7379 = w_sub02_result_dataout;
	assign w_sys_tmp7380 = (w_sys_tmp7381 + r_run_k_33);
	assign w_sys_tmp7381 = (r_run_copy0_j_163 * w_sys_tmp7378);
	assign w_sys_tmp7383 = (r_run_copy0_j_163 + w_sys_intOne);
	assign w_sys_tmp7384 = (r_run_copy1_j_164 + w_sys_intOne);
	assign w_sys_tmp7385 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp7464 = 32'sh00000031;
	assign w_sys_tmp7465 = ( !w_sys_tmp7466 );
	assign w_sys_tmp7466 = (w_sys_tmp7467 < r_run_j_34);
	assign w_sys_tmp7467 = 32'sh00000040;
	assign w_sys_tmp7469 = (r_run_j_34 - w_sys_tmp7470);
	assign w_sys_tmp7470 = 32'sh0000002f;
	assign w_sys_tmp7472 = (w_sys_tmp7473 + r_run_k_33);
	assign w_sys_tmp7473 = (r_run_copy1_j_166 * w_sys_tmp7474);
	assign w_sys_tmp7474 = 32'sh00000081;
	assign w_sys_tmp7475 = w_sub03_result_dataout;
	assign w_sys_tmp7476 = (w_sys_tmp7477 + r_run_k_33);
	assign w_sys_tmp7477 = (r_run_copy0_j_165 * w_sys_tmp7474);
	assign w_sys_tmp7479 = (r_run_copy0_j_165 + w_sys_intOne);
	assign w_sys_tmp7480 = (r_run_copy1_j_166 + w_sys_intOne);
	assign w_sys_tmp7481 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp7560 = 32'sh00000041;
	assign w_sys_tmp7561 = ( !w_sys_tmp7562 );
	assign w_sys_tmp7562 = (w_sys_tmp7563 < r_run_j_34);
	assign w_sys_tmp7563 = 32'sh00000050;
	assign w_sys_tmp7565 = (r_run_j_34 - w_sys_tmp7566);
	assign w_sys_tmp7566 = 32'sh0000003f;
	assign w_sys_tmp7568 = (w_sys_tmp7569 + r_run_k_33);
	assign w_sys_tmp7569 = (r_run_copy1_j_168 * w_sys_tmp7570);
	assign w_sys_tmp7570 = 32'sh00000081;
	assign w_sys_tmp7571 = w_sub04_result_dataout;
	assign w_sys_tmp7572 = (w_sys_tmp7573 + r_run_k_33);
	assign w_sys_tmp7573 = (r_run_copy0_j_167 * w_sys_tmp7570);
	assign w_sys_tmp7575 = (r_run_copy0_j_167 + w_sys_intOne);
	assign w_sys_tmp7576 = (r_run_copy1_j_168 + w_sys_intOne);
	assign w_sys_tmp7577 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp7656 = 32'sh00000051;
	assign w_sys_tmp7657 = ( !w_sys_tmp7658 );
	assign w_sys_tmp7658 = (w_sys_tmp7659 < r_run_j_34);
	assign w_sys_tmp7659 = 32'sh00000060;
	assign w_sys_tmp7661 = (r_run_j_34 - w_sys_tmp7662);
	assign w_sys_tmp7662 = 32'sh0000004f;
	assign w_sys_tmp7664 = (w_sys_tmp7665 + r_run_k_33);
	assign w_sys_tmp7665 = (r_run_copy1_j_170 * w_sys_tmp7666);
	assign w_sys_tmp7666 = 32'sh00000081;
	assign w_sys_tmp7667 = w_sub05_result_dataout;
	assign w_sys_tmp7668 = (w_sys_tmp7669 + r_run_k_33);
	assign w_sys_tmp7669 = (r_run_copy0_j_169 * w_sys_tmp7666);
	assign w_sys_tmp7671 = (r_run_copy0_j_169 + w_sys_intOne);
	assign w_sys_tmp7672 = (r_run_copy1_j_170 + w_sys_intOne);
	assign w_sys_tmp7673 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp7752 = 32'sh00000061;
	assign w_sys_tmp7753 = ( !w_sys_tmp7754 );
	assign w_sys_tmp7754 = (w_sys_tmp7755 < r_run_j_34);
	assign w_sys_tmp7755 = 32'sh00000070;
	assign w_sys_tmp7757 = (r_run_j_34 - w_sys_tmp7758);
	assign w_sys_tmp7758 = 32'sh0000005f;
	assign w_sys_tmp7760 = (w_sys_tmp7761 + r_run_k_33);
	assign w_sys_tmp7761 = (r_run_copy1_j_172 * w_sys_tmp7762);
	assign w_sys_tmp7762 = 32'sh00000081;
	assign w_sys_tmp7763 = w_sub06_result_dataout;
	assign w_sys_tmp7764 = (w_sys_tmp7765 + r_run_k_33);
	assign w_sys_tmp7765 = (r_run_copy0_j_171 * w_sys_tmp7762);
	assign w_sys_tmp7767 = (r_run_copy0_j_171 + w_sys_intOne);
	assign w_sys_tmp7768 = (r_run_copy1_j_172 + w_sys_intOne);
	assign w_sys_tmp7769 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp7848 = 32'sh00000071;
	assign w_sys_tmp7849 = ( !w_sys_tmp7850 );
	assign w_sys_tmp7850 = (w_sys_tmp7851 < r_run_j_34);
	assign w_sys_tmp7851 = 32'sh00000080;
	assign w_sys_tmp7853 = (r_run_j_34 - w_sys_tmp7854);
	assign w_sys_tmp7854 = 32'sh0000006f;
	assign w_sys_tmp7856 = (w_sys_tmp7857 + r_run_k_33);
	assign w_sys_tmp7857 = (r_run_copy1_j_174 * w_sys_tmp7858);
	assign w_sys_tmp7858 = 32'sh00000081;
	assign w_sys_tmp7859 = w_sub07_result_dataout;
	assign w_sys_tmp7860 = (w_sys_tmp7861 + r_run_k_33);
	assign w_sys_tmp7861 = (r_run_copy0_j_173 * w_sys_tmp7858);
	assign w_sys_tmp7863 = (r_run_copy0_j_173 + w_sys_intOne);
	assign w_sys_tmp7864 = (r_run_copy1_j_174 + w_sys_intOne);
	assign w_sys_tmp7865 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp7944 = 32'sh00000021;
	assign w_sys_tmp7945 = ( !w_sys_tmp7946 );
	assign w_sys_tmp7946 = (w_sys_tmp7947 < r_run_k_33);
	assign w_sys_tmp7947 = 32'sh00000040;
	assign w_sys_tmp7948 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp7949 = 32'sh00000002;
	assign w_sys_tmp7950 = ( !w_sys_tmp7951 );
	assign w_sys_tmp7951 = (w_sys_tmp7952 < r_run_j_34);
	assign w_sys_tmp7952 = 32'sh00000010;
	assign w_sys_tmp7955 = (w_sys_tmp7956 + r_run_k_33);
	assign w_sys_tmp7956 = (r_run_j_34 * w_sys_tmp7957);
	assign w_sys_tmp7957 = 32'sh00000081;
	assign w_sys_tmp7958 = w_sub08_result_dataout;
	assign w_sys_tmp7959 = (w_sys_tmp7960 + r_run_k_33);
	assign w_sys_tmp7960 = (r_run_copy0_j_175 * w_sys_tmp7957);
	assign w_sys_tmp7962 = (r_run_copy0_j_175 + w_sys_intOne);
	assign w_sys_tmp7963 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8024 = 32'sh00000011;
	assign w_sys_tmp8025 = ( !w_sys_tmp8026 );
	assign w_sys_tmp8026 = (w_sys_tmp8027 < r_run_j_34);
	assign w_sys_tmp8027 = 32'sh00000020;
	assign w_sys_tmp8029 = (r_run_j_34 - w_sys_tmp8030);
	assign w_sys_tmp8030 = 32'sh0000000f;
	assign w_sys_tmp8032 = (w_sys_tmp8033 + r_run_k_33);
	assign w_sys_tmp8033 = (r_run_copy1_j_177 * w_sys_tmp8034);
	assign w_sys_tmp8034 = 32'sh00000081;
	assign w_sys_tmp8035 = w_sub09_result_dataout;
	assign w_sys_tmp8036 = (w_sys_tmp8037 + r_run_k_33);
	assign w_sys_tmp8037 = (r_run_copy0_j_176 * w_sys_tmp8034);
	assign w_sys_tmp8039 = (r_run_copy0_j_176 + w_sys_intOne);
	assign w_sys_tmp8040 = (r_run_copy1_j_177 + w_sys_intOne);
	assign w_sys_tmp8041 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8120 = 32'sh00000021;
	assign w_sys_tmp8121 = ( !w_sys_tmp8122 );
	assign w_sys_tmp8122 = (w_sys_tmp8123 < r_run_j_34);
	assign w_sys_tmp8123 = 32'sh00000030;
	assign w_sys_tmp8125 = (r_run_j_34 - w_sys_tmp8126);
	assign w_sys_tmp8126 = 32'sh0000001f;
	assign w_sys_tmp8128 = (w_sys_tmp8129 + r_run_k_33);
	assign w_sys_tmp8129 = (r_run_copy1_j_179 * w_sys_tmp8130);
	assign w_sys_tmp8130 = 32'sh00000081;
	assign w_sys_tmp8131 = w_sub10_result_dataout;
	assign w_sys_tmp8132 = (w_sys_tmp8133 + r_run_k_33);
	assign w_sys_tmp8133 = (r_run_copy0_j_178 * w_sys_tmp8130);
	assign w_sys_tmp8135 = (r_run_copy0_j_178 + w_sys_intOne);
	assign w_sys_tmp8136 = (r_run_copy1_j_179 + w_sys_intOne);
	assign w_sys_tmp8137 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8216 = 32'sh00000031;
	assign w_sys_tmp8217 = ( !w_sys_tmp8218 );
	assign w_sys_tmp8218 = (w_sys_tmp8219 < r_run_j_34);
	assign w_sys_tmp8219 = 32'sh00000040;
	assign w_sys_tmp8221 = (r_run_j_34 - w_sys_tmp8222);
	assign w_sys_tmp8222 = 32'sh0000002f;
	assign w_sys_tmp8224 = (w_sys_tmp8225 + r_run_k_33);
	assign w_sys_tmp8225 = (r_run_copy1_j_181 * w_sys_tmp8226);
	assign w_sys_tmp8226 = 32'sh00000081;
	assign w_sys_tmp8227 = w_sub11_result_dataout;
	assign w_sys_tmp8228 = (w_sys_tmp8229 + r_run_k_33);
	assign w_sys_tmp8229 = (r_run_copy0_j_180 * w_sys_tmp8226);
	assign w_sys_tmp8231 = (r_run_copy0_j_180 + w_sys_intOne);
	assign w_sys_tmp8232 = (r_run_copy1_j_181 + w_sys_intOne);
	assign w_sys_tmp8233 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8312 = 32'sh00000041;
	assign w_sys_tmp8313 = ( !w_sys_tmp8314 );
	assign w_sys_tmp8314 = (w_sys_tmp8315 < r_run_j_34);
	assign w_sys_tmp8315 = 32'sh00000050;
	assign w_sys_tmp8317 = (r_run_j_34 - w_sys_tmp8318);
	assign w_sys_tmp8318 = 32'sh0000003f;
	assign w_sys_tmp8320 = (w_sys_tmp8321 + r_run_k_33);
	assign w_sys_tmp8321 = (r_run_copy1_j_183 * w_sys_tmp8322);
	assign w_sys_tmp8322 = 32'sh00000081;
	assign w_sys_tmp8323 = w_sub12_result_dataout;
	assign w_sys_tmp8324 = (w_sys_tmp8325 + r_run_k_33);
	assign w_sys_tmp8325 = (r_run_copy0_j_182 * w_sys_tmp8322);
	assign w_sys_tmp8327 = (r_run_copy0_j_182 + w_sys_intOne);
	assign w_sys_tmp8328 = (r_run_copy1_j_183 + w_sys_intOne);
	assign w_sys_tmp8329 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8408 = 32'sh00000051;
	assign w_sys_tmp8409 = ( !w_sys_tmp8410 );
	assign w_sys_tmp8410 = (w_sys_tmp8411 < r_run_j_34);
	assign w_sys_tmp8411 = 32'sh00000060;
	assign w_sys_tmp8413 = (r_run_j_34 - w_sys_tmp8414);
	assign w_sys_tmp8414 = 32'sh0000004f;
	assign w_sys_tmp8416 = (w_sys_tmp8417 + r_run_k_33);
	assign w_sys_tmp8417 = (r_run_copy1_j_185 * w_sys_tmp8418);
	assign w_sys_tmp8418 = 32'sh00000081;
	assign w_sys_tmp8419 = w_sub13_result_dataout;
	assign w_sys_tmp8420 = (w_sys_tmp8421 + r_run_k_33);
	assign w_sys_tmp8421 = (r_run_copy0_j_184 * w_sys_tmp8418);
	assign w_sys_tmp8423 = (r_run_copy0_j_184 + w_sys_intOne);
	assign w_sys_tmp8424 = (r_run_copy1_j_185 + w_sys_intOne);
	assign w_sys_tmp8425 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8504 = 32'sh00000061;
	assign w_sys_tmp8505 = ( !w_sys_tmp8506 );
	assign w_sys_tmp8506 = (w_sys_tmp8507 < r_run_j_34);
	assign w_sys_tmp8507 = 32'sh00000070;
	assign w_sys_tmp8509 = (r_run_j_34 - w_sys_tmp8510);
	assign w_sys_tmp8510 = 32'sh0000005f;
	assign w_sys_tmp8512 = (w_sys_tmp8513 + r_run_k_33);
	assign w_sys_tmp8513 = (r_run_copy1_j_187 * w_sys_tmp8514);
	assign w_sys_tmp8514 = 32'sh00000081;
	assign w_sys_tmp8515 = w_sub14_result_dataout;
	assign w_sys_tmp8516 = (w_sys_tmp8517 + r_run_k_33);
	assign w_sys_tmp8517 = (r_run_copy0_j_186 * w_sys_tmp8514);
	assign w_sys_tmp8519 = (r_run_copy0_j_186 + w_sys_intOne);
	assign w_sys_tmp8520 = (r_run_copy1_j_187 + w_sys_intOne);
	assign w_sys_tmp8521 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8600 = 32'sh00000071;
	assign w_sys_tmp8601 = ( !w_sys_tmp8602 );
	assign w_sys_tmp8602 = (w_sys_tmp8603 < r_run_j_34);
	assign w_sys_tmp8603 = 32'sh00000080;
	assign w_sys_tmp8605 = (r_run_j_34 - w_sys_tmp8606);
	assign w_sys_tmp8606 = 32'sh0000006f;
	assign w_sys_tmp8608 = (w_sys_tmp8609 + r_run_k_33);
	assign w_sys_tmp8609 = (r_run_copy1_j_189 * w_sys_tmp8610);
	assign w_sys_tmp8610 = 32'sh00000081;
	assign w_sys_tmp8611 = w_sub15_result_dataout;
	assign w_sys_tmp8612 = (w_sys_tmp8613 + r_run_k_33);
	assign w_sys_tmp8613 = (r_run_copy0_j_188 * w_sys_tmp8610);
	assign w_sys_tmp8615 = (r_run_copy0_j_188 + w_sys_intOne);
	assign w_sys_tmp8616 = (r_run_copy1_j_189 + w_sys_intOne);
	assign w_sys_tmp8617 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8696 = 32'sh00000041;
	assign w_sys_tmp8697 = ( !w_sys_tmp8698 );
	assign w_sys_tmp8698 = (w_sys_tmp8699 < r_run_k_33);
	assign w_sys_tmp8699 = 32'sh00000060;
	assign w_sys_tmp8700 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp8701 = 32'sh00000002;
	assign w_sys_tmp8702 = ( !w_sys_tmp8703 );
	assign w_sys_tmp8703 = (w_sys_tmp8704 < r_run_j_34);
	assign w_sys_tmp8704 = 32'sh00000010;
	assign w_sys_tmp8707 = (w_sys_tmp8708 + r_run_k_33);
	assign w_sys_tmp8708 = (r_run_j_34 * w_sys_tmp8709);
	assign w_sys_tmp8709 = 32'sh00000081;
	assign w_sys_tmp8710 = w_sub16_result_dataout;
	assign w_sys_tmp8711 = (w_sys_tmp8712 + r_run_k_33);
	assign w_sys_tmp8712 = (r_run_copy0_j_190 * w_sys_tmp8709);
	assign w_sys_tmp8714 = (r_run_copy0_j_190 + w_sys_intOne);
	assign w_sys_tmp8715 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8776 = 32'sh00000011;
	assign w_sys_tmp8777 = ( !w_sys_tmp8778 );
	assign w_sys_tmp8778 = (w_sys_tmp8779 < r_run_j_34);
	assign w_sys_tmp8779 = 32'sh00000020;
	assign w_sys_tmp8781 = (r_run_j_34 - w_sys_tmp8782);
	assign w_sys_tmp8782 = 32'sh0000000f;
	assign w_sys_tmp8784 = (w_sys_tmp8785 + r_run_k_33);
	assign w_sys_tmp8785 = (r_run_copy1_j_192 * w_sys_tmp8786);
	assign w_sys_tmp8786 = 32'sh00000081;
	assign w_sys_tmp8787 = w_sub17_result_dataout;
	assign w_sys_tmp8788 = (w_sys_tmp8789 + r_run_k_33);
	assign w_sys_tmp8789 = (r_run_copy0_j_191 * w_sys_tmp8786);
	assign w_sys_tmp8791 = (r_run_copy0_j_191 + w_sys_intOne);
	assign w_sys_tmp8792 = (r_run_copy1_j_192 + w_sys_intOne);
	assign w_sys_tmp8793 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8872 = 32'sh00000021;
	assign w_sys_tmp8873 = ( !w_sys_tmp8874 );
	assign w_sys_tmp8874 = (w_sys_tmp8875 < r_run_j_34);
	assign w_sys_tmp8875 = 32'sh00000030;
	assign w_sys_tmp8877 = (r_run_j_34 - w_sys_tmp8878);
	assign w_sys_tmp8878 = 32'sh0000001f;
	assign w_sys_tmp8880 = (w_sys_tmp8881 + r_run_k_33);
	assign w_sys_tmp8881 = (r_run_copy1_j_194 * w_sys_tmp8882);
	assign w_sys_tmp8882 = 32'sh00000081;
	assign w_sys_tmp8883 = w_sub18_result_dataout;
	assign w_sys_tmp8884 = (w_sys_tmp8885 + r_run_k_33);
	assign w_sys_tmp8885 = (r_run_copy0_j_193 * w_sys_tmp8882);
	assign w_sys_tmp8887 = (r_run_copy0_j_193 + w_sys_intOne);
	assign w_sys_tmp8888 = (r_run_copy1_j_194 + w_sys_intOne);
	assign w_sys_tmp8889 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp8968 = 32'sh00000031;
	assign w_sys_tmp8969 = ( !w_sys_tmp8970 );
	assign w_sys_tmp8970 = (w_sys_tmp8971 < r_run_j_34);
	assign w_sys_tmp8971 = 32'sh00000040;
	assign w_sys_tmp8973 = (r_run_j_34 - w_sys_tmp8974);
	assign w_sys_tmp8974 = 32'sh0000002f;
	assign w_sys_tmp8976 = (w_sys_tmp8977 + r_run_k_33);
	assign w_sys_tmp8977 = (r_run_copy1_j_196 * w_sys_tmp8978);
	assign w_sys_tmp8978 = 32'sh00000081;
	assign w_sys_tmp8979 = w_sub19_result_dataout;
	assign w_sys_tmp8980 = (w_sys_tmp8981 + r_run_k_33);
	assign w_sys_tmp8981 = (r_run_copy0_j_195 * w_sys_tmp8978);
	assign w_sys_tmp8983 = (r_run_copy0_j_195 + w_sys_intOne);
	assign w_sys_tmp8984 = (r_run_copy1_j_196 + w_sys_intOne);
	assign w_sys_tmp8985 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp9064 = 32'sh00000041;
	assign w_sys_tmp9065 = ( !w_sys_tmp9066 );
	assign w_sys_tmp9066 = (w_sys_tmp9067 < r_run_j_34);
	assign w_sys_tmp9067 = 32'sh00000050;
	assign w_sys_tmp9069 = (r_run_j_34 - w_sys_tmp9070);
	assign w_sys_tmp9070 = 32'sh0000003f;
	assign w_sys_tmp9072 = (w_sys_tmp9073 + r_run_k_33);
	assign w_sys_tmp9073 = (r_run_copy1_j_198 * w_sys_tmp9074);
	assign w_sys_tmp9074 = 32'sh00000081;
	assign w_sys_tmp9075 = w_sub20_result_dataout;
	assign w_sys_tmp9076 = (w_sys_tmp9077 + r_run_k_33);
	assign w_sys_tmp9077 = (r_run_copy0_j_197 * w_sys_tmp9074);
	assign w_sys_tmp9079 = (r_run_copy0_j_197 + w_sys_intOne);
	assign w_sys_tmp9080 = (r_run_copy1_j_198 + w_sys_intOne);
	assign w_sys_tmp9081 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp9160 = 32'sh00000051;
	assign w_sys_tmp9161 = ( !w_sys_tmp9162 );
	assign w_sys_tmp9162 = (w_sys_tmp9163 < r_run_j_34);
	assign w_sys_tmp9163 = 32'sh00000060;
	assign w_sys_tmp9165 = (r_run_j_34 - w_sys_tmp9166);
	assign w_sys_tmp9166 = 32'sh0000004f;
	assign w_sys_tmp9168 = (w_sys_tmp9169 + r_run_k_33);
	assign w_sys_tmp9169 = (r_run_copy1_j_200 * w_sys_tmp9170);
	assign w_sys_tmp9170 = 32'sh00000081;
	assign w_sys_tmp9171 = w_sub21_result_dataout;
	assign w_sys_tmp9172 = (w_sys_tmp9173 + r_run_k_33);
	assign w_sys_tmp9173 = (r_run_copy0_j_199 * w_sys_tmp9170);
	assign w_sys_tmp9175 = (r_run_copy0_j_199 + w_sys_intOne);
	assign w_sys_tmp9176 = (r_run_copy1_j_200 + w_sys_intOne);
	assign w_sys_tmp9177 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp9256 = 32'sh00000061;
	assign w_sys_tmp9257 = ( !w_sys_tmp9258 );
	assign w_sys_tmp9258 = (w_sys_tmp9259 < r_run_j_34);
	assign w_sys_tmp9259 = 32'sh00000070;
	assign w_sys_tmp9261 = (r_run_j_34 - w_sys_tmp9262);
	assign w_sys_tmp9262 = 32'sh0000005f;
	assign w_sys_tmp9264 = (w_sys_tmp9265 + r_run_k_33);
	assign w_sys_tmp9265 = (r_run_copy1_j_202 * w_sys_tmp9266);
	assign w_sys_tmp9266 = 32'sh00000081;
	assign w_sys_tmp9267 = w_sub22_result_dataout;
	assign w_sys_tmp9268 = (w_sys_tmp9269 + r_run_k_33);
	assign w_sys_tmp9269 = (r_run_copy0_j_201 * w_sys_tmp9266);
	assign w_sys_tmp9271 = (r_run_copy0_j_201 + w_sys_intOne);
	assign w_sys_tmp9272 = (r_run_copy1_j_202 + w_sys_intOne);
	assign w_sys_tmp9273 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp9352 = 32'sh00000071;
	assign w_sys_tmp9353 = ( !w_sys_tmp9354 );
	assign w_sys_tmp9354 = (w_sys_tmp9355 < r_run_j_34);
	assign w_sys_tmp9355 = 32'sh00000080;
	assign w_sys_tmp9357 = (r_run_j_34 - w_sys_tmp9358);
	assign w_sys_tmp9358 = 32'sh0000006f;
	assign w_sys_tmp9360 = (w_sys_tmp9361 + r_run_k_33);
	assign w_sys_tmp9361 = (r_run_copy1_j_204 * w_sys_tmp9362);
	assign w_sys_tmp9362 = 32'sh00000081;
	assign w_sys_tmp9363 = w_sub23_result_dataout;
	assign w_sys_tmp9364 = (w_sys_tmp9365 + r_run_k_33);
	assign w_sys_tmp9365 = (r_run_copy0_j_203 * w_sys_tmp9362);
	assign w_sys_tmp9367 = (r_run_copy0_j_203 + w_sys_intOne);
	assign w_sys_tmp9368 = (r_run_copy1_j_204 + w_sys_intOne);
	assign w_sys_tmp9369 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp9448 = 32'sh00000061;
	assign w_sys_tmp9449 = ( !w_sys_tmp9450 );
	assign w_sys_tmp9450 = (w_sys_tmp9451 < r_run_k_33);
	assign w_sys_tmp9451 = 32'sh00000080;
	assign w_sys_tmp9452 = (r_run_k_33 + w_sys_intOne);
	assign w_sys_tmp9453 = 32'sh00000002;
	assign w_sys_tmp9454 = ( !w_sys_tmp9455 );
	assign w_sys_tmp9455 = (w_sys_tmp9456 < r_run_j_34);
	assign w_sys_tmp9456 = 32'sh00000010;
	assign w_sys_tmp9459 = (w_sys_tmp9460 + r_run_k_33);
	assign w_sys_tmp9460 = (r_run_j_34 * w_sys_tmp9461);
	assign w_sys_tmp9461 = 32'sh00000081;
	assign w_sys_tmp9462 = w_sub24_result_dataout;
	assign w_sys_tmp9463 = (w_sys_tmp9464 + r_run_k_33);
	assign w_sys_tmp9464 = (r_run_copy0_j_205 * w_sys_tmp9461);
	assign w_sys_tmp9466 = (r_run_copy0_j_205 + w_sys_intOne);
	assign w_sys_tmp9467 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp9528 = 32'sh00000011;
	assign w_sys_tmp9529 = ( !w_sys_tmp9530 );
	assign w_sys_tmp9530 = (w_sys_tmp9531 < r_run_j_34);
	assign w_sys_tmp9531 = 32'sh00000020;
	assign w_sys_tmp9533 = (r_run_j_34 - w_sys_tmp9534);
	assign w_sys_tmp9534 = 32'sh0000000f;
	assign w_sys_tmp9536 = (w_sys_tmp9537 + r_run_k_33);
	assign w_sys_tmp9537 = (r_run_copy1_j_207 * w_sys_tmp9538);
	assign w_sys_tmp9538 = 32'sh00000081;
	assign w_sys_tmp9539 = w_sub25_result_dataout;
	assign w_sys_tmp9540 = (w_sys_tmp9541 + r_run_k_33);
	assign w_sys_tmp9541 = (r_run_copy0_j_206 * w_sys_tmp9538);
	assign w_sys_tmp9543 = (r_run_copy0_j_206 + w_sys_intOne);
	assign w_sys_tmp9544 = (r_run_copy1_j_207 + w_sys_intOne);
	assign w_sys_tmp9545 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp9624 = 32'sh00000021;
	assign w_sys_tmp9625 = ( !w_sys_tmp9626 );
	assign w_sys_tmp9626 = (w_sys_tmp9627 < r_run_j_34);
	assign w_sys_tmp9627 = 32'sh00000030;
	assign w_sys_tmp9629 = (r_run_j_34 - w_sys_tmp9630);
	assign w_sys_tmp9630 = 32'sh0000001f;
	assign w_sys_tmp9632 = (w_sys_tmp9633 + r_run_k_33);
	assign w_sys_tmp9633 = (r_run_copy1_j_209 * w_sys_tmp9634);
	assign w_sys_tmp9634 = 32'sh00000081;
	assign w_sys_tmp9635 = w_sub26_result_dataout;
	assign w_sys_tmp9636 = (w_sys_tmp9637 + r_run_k_33);
	assign w_sys_tmp9637 = (r_run_copy0_j_208 * w_sys_tmp9634);
	assign w_sys_tmp9639 = (r_run_copy0_j_208 + w_sys_intOne);
	assign w_sys_tmp9640 = (r_run_copy1_j_209 + w_sys_intOne);
	assign w_sys_tmp9641 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp9720 = 32'sh00000031;
	assign w_sys_tmp9721 = ( !w_sys_tmp9722 );
	assign w_sys_tmp9722 = (w_sys_tmp9723 < r_run_j_34);
	assign w_sys_tmp9723 = 32'sh00000040;
	assign w_sys_tmp9725 = (r_run_j_34 - w_sys_tmp9726);
	assign w_sys_tmp9726 = 32'sh0000002f;
	assign w_sys_tmp9728 = (w_sys_tmp9729 + r_run_k_33);
	assign w_sys_tmp9729 = (r_run_copy1_j_211 * w_sys_tmp9730);
	assign w_sys_tmp9730 = 32'sh00000081;
	assign w_sys_tmp9731 = w_sub27_result_dataout;
	assign w_sys_tmp9732 = (w_sys_tmp9733 + r_run_k_33);
	assign w_sys_tmp9733 = (r_run_copy0_j_210 * w_sys_tmp9730);
	assign w_sys_tmp9735 = (r_run_copy0_j_210 + w_sys_intOne);
	assign w_sys_tmp9736 = (r_run_copy1_j_211 + w_sys_intOne);
	assign w_sys_tmp9737 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp9816 = 32'sh00000041;
	assign w_sys_tmp9817 = ( !w_sys_tmp9818 );
	assign w_sys_tmp9818 = (w_sys_tmp9819 < r_run_j_34);
	assign w_sys_tmp9819 = 32'sh00000050;
	assign w_sys_tmp9821 = (r_run_j_34 - w_sys_tmp9822);
	assign w_sys_tmp9822 = 32'sh0000003f;
	assign w_sys_tmp9824 = (w_sys_tmp9825 + r_run_k_33);
	assign w_sys_tmp9825 = (r_run_copy1_j_213 * w_sys_tmp9826);
	assign w_sys_tmp9826 = 32'sh00000081;
	assign w_sys_tmp9827 = w_sub28_result_dataout;
	assign w_sys_tmp9828 = (w_sys_tmp9829 + r_run_k_33);
	assign w_sys_tmp9829 = (r_run_copy0_j_212 * w_sys_tmp9826);
	assign w_sys_tmp9831 = (r_run_copy0_j_212 + w_sys_intOne);
	assign w_sys_tmp9832 = (r_run_copy1_j_213 + w_sys_intOne);
	assign w_sys_tmp9833 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp9912 = 32'sh00000051;
	assign w_sys_tmp9913 = ( !w_sys_tmp9914 );
	assign w_sys_tmp9914 = (w_sys_tmp9915 < r_run_j_34);
	assign w_sys_tmp9915 = 32'sh00000060;
	assign w_sys_tmp9917 = (r_run_j_34 - w_sys_tmp9918);
	assign w_sys_tmp9918 = 32'sh0000004f;
	assign w_sys_tmp9920 = (w_sys_tmp9921 + r_run_k_33);
	assign w_sys_tmp9921 = (r_run_copy1_j_215 * w_sys_tmp9922);
	assign w_sys_tmp9922 = 32'sh00000081;
	assign w_sys_tmp9923 = w_sub29_result_dataout;
	assign w_sys_tmp9924 = (w_sys_tmp9925 + r_run_k_33);
	assign w_sys_tmp9925 = (r_run_copy0_j_214 * w_sys_tmp9922);
	assign w_sys_tmp9927 = (r_run_copy0_j_214 + w_sys_intOne);
	assign w_sys_tmp9928 = (r_run_copy1_j_215 + w_sys_intOne);
	assign w_sys_tmp9929 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp10008 = 32'sh00000061;
	assign w_sys_tmp10009 = ( !w_sys_tmp10010 );
	assign w_sys_tmp10010 = (w_sys_tmp10011 < r_run_j_34);
	assign w_sys_tmp10011 = 32'sh00000070;
	assign w_sys_tmp10013 = (r_run_j_34 - w_sys_tmp10014);
	assign w_sys_tmp10014 = 32'sh0000005f;
	assign w_sys_tmp10016 = (w_sys_tmp10017 + r_run_k_33);
	assign w_sys_tmp10017 = (r_run_copy1_j_217 * w_sys_tmp10018);
	assign w_sys_tmp10018 = 32'sh00000081;
	assign w_sys_tmp10019 = w_sub30_result_dataout;
	assign w_sys_tmp10020 = (w_sys_tmp10021 + r_run_k_33);
	assign w_sys_tmp10021 = (r_run_copy0_j_216 * w_sys_tmp10018);
	assign w_sys_tmp10023 = (r_run_copy0_j_216 + w_sys_intOne);
	assign w_sys_tmp10024 = (r_run_copy1_j_217 + w_sys_intOne);
	assign w_sys_tmp10025 = (r_run_j_34 + w_sys_intOne);
	assign w_sys_tmp10104 = 32'sh00000071;
	assign w_sys_tmp10105 = ( !w_sys_tmp10106 );
	assign w_sys_tmp10106 = (w_sys_tmp10107 < r_run_j_34);
	assign w_sys_tmp10107 = 32'sh00000080;
	assign w_sys_tmp10109 = (r_run_j_34 - w_sys_tmp10110);
	assign w_sys_tmp10110 = 32'sh0000006f;
	assign w_sys_tmp10112 = (w_sys_tmp10113 + r_run_k_33);
	assign w_sys_tmp10113 = (r_run_copy1_j_219 * w_sys_tmp10114);
	assign w_sys_tmp10114 = 32'sh00000081;
	assign w_sys_tmp10115 = w_sub31_result_dataout;
	assign w_sys_tmp10116 = (w_sys_tmp10117 + r_run_k_33);
	assign w_sys_tmp10117 = (r_run_copy0_j_218 * w_sys_tmp10114);
	assign w_sys_tmp10119 = (r_run_copy0_j_218 + w_sys_intOne);
	assign w_sys_tmp10120 = (r_run_copy1_j_219 + w_sys_intOne);
	assign w_sys_tmp10121 = (r_run_j_34 + w_sys_intOne);


	sub19
		sub19_inst(
			.i_fld_result_1_addr_0 (w_sub19_result_addr),
			.i_fld_result_1_datain_0 (w_sub19_result_datain),
			.o_fld_result_1_dataout_0 (w_sub19_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub19_result_r_w),
			.i_fld_u_0_addr_0 (w_sub19_u_addr),
			.i_fld_u_0_datain_0 (w_sub19_u_datain),
			.o_fld_u_0_dataout_0 (w_sub19_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub19_u_r_w),
			.o_run_busy (w_sub19_run_busy),
			.i_run_req (r_sub19_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_result_1_addr_0 (w_sub12_result_addr),
			.i_fld_result_1_datain_0 (w_sub12_result_datain),
			.o_fld_result_1_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub12_result_r_w),
			.i_fld_u_0_addr_0 (w_sub12_u_addr),
			.i_fld_u_0_datain_0 (w_sub12_u_datain),
			.o_fld_u_0_dataout_0 (w_sub12_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub12_u_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_result_1_addr_0 (w_sub11_result_addr),
			.i_fld_result_1_datain_0 (w_sub11_result_datain),
			.o_fld_result_1_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub11_result_r_w),
			.i_fld_u_0_addr_0 (w_sub11_u_addr),
			.i_fld_u_0_datain_0 (w_sub11_u_datain),
			.o_fld_u_0_dataout_0 (w_sub11_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub11_u_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_result_1_addr_0 (w_sub14_result_addr),
			.i_fld_result_1_datain_0 (w_sub14_result_datain),
			.o_fld_result_1_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub14_result_r_w),
			.i_fld_u_0_addr_0 (w_sub14_u_addr),
			.i_fld_u_0_datain_0 (w_sub14_u_datain),
			.o_fld_u_0_dataout_0 (w_sub14_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub14_u_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_result_1_addr_0 (w_sub13_result_addr),
			.i_fld_result_1_datain_0 (w_sub13_result_datain),
			.o_fld_result_1_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub13_result_r_w),
			.i_fld_u_0_addr_0 (w_sub13_u_addr),
			.i_fld_u_0_datain_0 (w_sub13_u_datain),
			.o_fld_u_0_dataout_0 (w_sub13_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub13_u_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub16
		sub16_inst(
			.i_fld_result_1_addr_0 (w_sub16_result_addr),
			.i_fld_result_1_datain_0 (w_sub16_result_datain),
			.o_fld_result_1_dataout_0 (w_sub16_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub16_result_r_w),
			.i_fld_u_0_addr_0 (w_sub16_u_addr),
			.i_fld_u_0_datain_0 (w_sub16_u_datain),
			.o_fld_u_0_dataout_0 (w_sub16_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub16_u_r_w),
			.o_run_busy (w_sub16_run_busy),
			.i_run_req (r_sub16_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_result_1_addr_0 (w_sub15_result_addr),
			.i_fld_result_1_datain_0 (w_sub15_result_datain),
			.o_fld_result_1_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub15_result_r_w),
			.i_fld_u_0_addr_0 (w_sub15_u_addr),
			.i_fld_u_0_datain_0 (w_sub15_u_datain),
			.o_fld_u_0_dataout_0 (w_sub15_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub15_u_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub18
		sub18_inst(
			.i_fld_result_1_addr_0 (w_sub18_result_addr),
			.i_fld_result_1_datain_0 (w_sub18_result_datain),
			.o_fld_result_1_dataout_0 (w_sub18_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub18_result_r_w),
			.i_fld_u_0_addr_0 (w_sub18_u_addr),
			.i_fld_u_0_datain_0 (w_sub18_u_datain),
			.o_fld_u_0_dataout_0 (w_sub18_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub18_u_r_w),
			.o_run_busy (w_sub18_run_busy),
			.i_run_req (r_sub18_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub17
		sub17_inst(
			.i_fld_result_1_addr_0 (w_sub17_result_addr),
			.i_fld_result_1_datain_0 (w_sub17_result_datain),
			.o_fld_result_1_dataout_0 (w_sub17_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub17_result_r_w),
			.i_fld_u_0_addr_0 (w_sub17_u_addr),
			.i_fld_u_0_datain_0 (w_sub17_u_datain),
			.o_fld_u_0_dataout_0 (w_sub17_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub17_u_r_w),
			.o_run_busy (w_sub17_run_busy),
			.i_run_req (r_sub17_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub20
		sub20_inst(
			.i_fld_result_1_addr_0 (w_sub20_result_addr),
			.i_fld_result_1_datain_0 (w_sub20_result_datain),
			.o_fld_result_1_dataout_0 (w_sub20_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub20_result_r_w),
			.i_fld_u_0_addr_0 (w_sub20_u_addr),
			.i_fld_u_0_datain_0 (w_sub20_u_datain),
			.o_fld_u_0_dataout_0 (w_sub20_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub20_u_r_w),
			.o_run_busy (w_sub20_run_busy),
			.i_run_req (r_sub20_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub21
		sub21_inst(
			.i_fld_result_1_addr_0 (w_sub21_result_addr),
			.i_fld_result_1_datain_0 (w_sub21_result_datain),
			.o_fld_result_1_dataout_0 (w_sub21_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub21_result_r_w),
			.i_fld_u_0_addr_0 (w_sub21_u_addr),
			.i_fld_u_0_datain_0 (w_sub21_u_datain),
			.o_fld_u_0_dataout_0 (w_sub21_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub21_u_r_w),
			.o_run_busy (w_sub21_run_busy),
			.i_run_req (r_sub21_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub28
		sub28_inst(
			.i_fld_result_1_addr_0 (w_sub28_result_addr),
			.i_fld_result_1_datain_0 (w_sub28_result_datain),
			.o_fld_result_1_dataout_0 (w_sub28_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub28_result_r_w),
			.i_fld_u_0_addr_0 (w_sub28_u_addr),
			.i_fld_u_0_datain_0 (w_sub28_u_datain),
			.o_fld_u_0_dataout_0 (w_sub28_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub28_u_r_w),
			.o_run_busy (w_sub28_run_busy),
			.i_run_req (r_sub28_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub29
		sub29_inst(
			.i_fld_result_1_addr_0 (w_sub29_result_addr),
			.i_fld_result_1_datain_0 (w_sub29_result_datain),
			.o_fld_result_1_dataout_0 (w_sub29_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub29_result_r_w),
			.i_fld_u_0_addr_0 (w_sub29_u_addr),
			.i_fld_u_0_datain_0 (w_sub29_u_datain),
			.o_fld_u_0_dataout_0 (w_sub29_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub29_u_r_w),
			.o_run_busy (w_sub29_run_busy),
			.i_run_req (r_sub29_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub26
		sub26_inst(
			.i_fld_result_1_addr_0 (w_sub26_result_addr),
			.i_fld_result_1_datain_0 (w_sub26_result_datain),
			.o_fld_result_1_dataout_0 (w_sub26_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub26_result_r_w),
			.i_fld_u_0_addr_0 (w_sub26_u_addr),
			.i_fld_u_0_datain_0 (w_sub26_u_datain),
			.o_fld_u_0_dataout_0 (w_sub26_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub26_u_r_w),
			.o_run_busy (w_sub26_run_busy),
			.i_run_req (r_sub26_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub09
		sub09_inst(
			.i_fld_result_1_addr_0 (w_sub09_result_addr),
			.i_fld_result_1_datain_0 (w_sub09_result_datain),
			.o_fld_result_1_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub09_result_r_w),
			.i_fld_u_0_addr_0 (w_sub09_u_addr),
			.i_fld_u_0_datain_0 (w_sub09_u_datain),
			.o_fld_u_0_dataout_0 (w_sub09_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub09_u_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub27
		sub27_inst(
			.i_fld_result_1_addr_0 (w_sub27_result_addr),
			.i_fld_result_1_datain_0 (w_sub27_result_datain),
			.o_fld_result_1_dataout_0 (w_sub27_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub27_result_r_w),
			.i_fld_u_0_addr_0 (w_sub27_u_addr),
			.i_fld_u_0_datain_0 (w_sub27_u_datain),
			.o_fld_u_0_dataout_0 (w_sub27_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub27_u_r_w),
			.o_run_busy (w_sub27_run_busy),
			.i_run_req (r_sub27_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_result_1_addr_0 (w_sub08_result_addr),
			.i_fld_result_1_datain_0 (w_sub08_result_datain),
			.o_fld_result_1_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub08_result_r_w),
			.i_fld_u_0_addr_0 (w_sub08_u_addr),
			.i_fld_u_0_datain_0 (w_sub08_u_datain),
			.o_fld_u_0_dataout_0 (w_sub08_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub08_u_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub24
		sub24_inst(
			.i_fld_result_1_addr_0 (w_sub24_result_addr),
			.i_fld_result_1_datain_0 (w_sub24_result_datain),
			.o_fld_result_1_dataout_0 (w_sub24_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub24_result_r_w),
			.i_fld_u_0_addr_0 (w_sub24_u_addr),
			.i_fld_u_0_datain_0 (w_sub24_u_datain),
			.o_fld_u_0_dataout_0 (w_sub24_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub24_u_r_w),
			.o_run_busy (w_sub24_run_busy),
			.i_run_req (r_sub24_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub25
		sub25_inst(
			.i_fld_result_1_addr_0 (w_sub25_result_addr),
			.i_fld_result_1_datain_0 (w_sub25_result_datain),
			.o_fld_result_1_dataout_0 (w_sub25_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub25_result_r_w),
			.i_fld_u_0_addr_0 (w_sub25_u_addr),
			.i_fld_u_0_datain_0 (w_sub25_u_datain),
			.o_fld_u_0_dataout_0 (w_sub25_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub25_u_r_w),
			.o_run_busy (w_sub25_run_busy),
			.i_run_req (r_sub25_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub22
		sub22_inst(
			.i_fld_result_1_addr_0 (w_sub22_result_addr),
			.i_fld_result_1_datain_0 (w_sub22_result_datain),
			.o_fld_result_1_dataout_0 (w_sub22_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub22_result_r_w),
			.i_fld_u_0_addr_0 (w_sub22_u_addr),
			.i_fld_u_0_datain_0 (w_sub22_u_datain),
			.o_fld_u_0_dataout_0 (w_sub22_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub22_u_r_w),
			.o_run_busy (w_sub22_run_busy),
			.i_run_req (r_sub22_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub23
		sub23_inst(
			.i_fld_result_1_addr_0 (w_sub23_result_addr),
			.i_fld_result_1_datain_0 (w_sub23_result_datain),
			.o_fld_result_1_dataout_0 (w_sub23_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub23_result_r_w),
			.i_fld_u_0_addr_0 (w_sub23_u_addr),
			.i_fld_u_0_datain_0 (w_sub23_u_datain),
			.o_fld_u_0_dataout_0 (w_sub23_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub23_u_r_w),
			.o_run_busy (w_sub23_run_busy),
			.i_run_req (r_sub23_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_result_1_addr_0 (w_sub03_result_addr),
			.i_fld_result_1_datain_0 (w_sub03_result_datain),
			.o_fld_result_1_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub03_result_r_w),
			.i_fld_u_0_addr_0 (w_sub03_u_addr),
			.i_fld_u_0_datain_0 (w_sub03_u_datain),
			.o_fld_u_0_dataout_0 (w_sub03_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub03_u_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_result_1_addr_0 (w_sub02_result_addr),
			.i_fld_result_1_datain_0 (w_sub02_result_datain),
			.o_fld_result_1_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub02_result_r_w),
			.i_fld_u_0_addr_0 (w_sub02_u_addr),
			.i_fld_u_0_datain_0 (w_sub02_u_datain),
			.o_fld_u_0_dataout_0 (w_sub02_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub02_u_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_result_1_addr_0 (w_sub01_result_addr),
			.i_fld_result_1_datain_0 (w_sub01_result_datain),
			.o_fld_result_1_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub01_result_r_w),
			.i_fld_u_0_addr_0 (w_sub01_u_addr),
			.i_fld_u_0_datain_0 (w_sub01_u_datain),
			.o_fld_u_0_dataout_0 (w_sub01_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub01_u_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_result_1_addr_0 (w_sub00_result_addr),
			.i_fld_result_1_datain_0 (w_sub00_result_datain),
			.o_fld_result_1_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub00_result_r_w),
			.i_fld_u_0_addr_0 (w_sub00_u_addr),
			.i_fld_u_0_datain_0 (w_sub00_u_datain),
			.o_fld_u_0_dataout_0 (w_sub00_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub00_u_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_result_1_addr_0 (w_sub07_result_addr),
			.i_fld_result_1_datain_0 (w_sub07_result_datain),
			.o_fld_result_1_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub07_result_r_w),
			.i_fld_u_0_addr_0 (w_sub07_u_addr),
			.i_fld_u_0_datain_0 (w_sub07_u_datain),
			.o_fld_u_0_dataout_0 (w_sub07_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub07_u_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_result_1_addr_0 (w_sub06_result_addr),
			.i_fld_result_1_datain_0 (w_sub06_result_datain),
			.o_fld_result_1_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub06_result_r_w),
			.i_fld_u_0_addr_0 (w_sub06_u_addr),
			.i_fld_u_0_datain_0 (w_sub06_u_datain),
			.o_fld_u_0_dataout_0 (w_sub06_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub06_u_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_result_1_addr_0 (w_sub05_result_addr),
			.i_fld_result_1_datain_0 (w_sub05_result_datain),
			.o_fld_result_1_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub05_result_r_w),
			.i_fld_u_0_addr_0 (w_sub05_u_addr),
			.i_fld_u_0_datain_0 (w_sub05_u_datain),
			.o_fld_u_0_dataout_0 (w_sub05_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub05_u_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_result_1_addr_0 (w_sub04_result_addr),
			.i_fld_result_1_datain_0 (w_sub04_result_datain),
			.o_fld_result_1_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub04_result_r_w),
			.i_fld_u_0_addr_0 (w_sub04_u_addr),
			.i_fld_u_0_datain_0 (w_sub04_u_datain),
			.o_fld_u_0_dataout_0 (w_sub04_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub04_u_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_result_1_addr_0 (w_sub10_result_addr),
			.i_fld_result_1_datain_0 (w_sub10_result_datain),
			.o_fld_result_1_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub10_result_r_w),
			.i_fld_u_0_addr_0 (w_sub10_u_addr),
			.i_fld_u_0_datain_0 (w_sub10_u_datain),
			.o_fld_u_0_dataout_0 (w_sub10_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub10_u_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub31
		sub31_inst(
			.i_fld_result_1_addr_0 (w_sub31_result_addr),
			.i_fld_result_1_datain_0 (w_sub31_result_datain),
			.o_fld_result_1_dataout_0 (w_sub31_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub31_result_r_w),
			.i_fld_u_0_addr_0 (w_sub31_u_addr),
			.i_fld_u_0_datain_0 (w_sub31_u_datain),
			.o_fld_u_0_dataout_0 (w_sub31_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub31_u_r_w),
			.o_run_busy (w_sub31_run_busy),
			.i_run_req (r_sub31_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub30
		sub30_inst(
			.i_fld_result_1_addr_0 (w_sub30_result_addr),
			.i_fld_result_1_datain_0 (w_sub30_result_datain),
			.o_fld_result_1_dataout_0 (w_sub30_result_dataout),
			.i_fld_result_1_r_w_0 (w_sub30_result_r_w),
			.i_fld_u_0_addr_0 (w_sub30_u_addr),
			.i_fld_u_0_datain_0 (w_sub30_u_datain),
			.o_fld_u_0_dataout_0 (w_sub30_u_dataout),
			.i_fld_u_0_r_w_0 (w_sub30_u_r_w),
			.o_run_busy (w_sub30_run_busy),
			.i_run_req (r_sub30_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(15), .WORDS(16900) )
		dpram_u_0(
			.clk (clock),
			.ce_0 (w_fld_u_0_ce_0),
			.addr_0 (w_fld_u_0_addr_0),
			.datain_0 (w_fld_u_0_datain_0),
			.dataout_0 (w_fld_u_0_dataout_0),
			.r_w_0 (w_fld_u_0_r_w_0),
			.ce_1 (w_fld_u_0_ce_1),
			.addr_1 (r_fld_u_0_addr_1),
			.datain_1 (r_fld_u_0_datain_1),
			.dataout_1 (w_fld_u_0_dataout_1),
			.r_w_1 (r_fld_u_0_r_w_1)
		);

	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						10'h207: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 10'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h0: begin
							r_sys_run_phase <= 10'h2;
						end

						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h4;

									end
								end

							endcase
						end

						10'h4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h5;

									end
								end

							endcase
						end

						10'h5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3) ? 10'h9 : 10'hf);

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h5;

									end
								end

							endcase
						end

						10'h9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'ha;

									end
								end

							endcase
						end

						10'ha: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6) ? 10'hd : 10'h6);

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_phase <= 10'ha;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h10;

									end
								end

							endcase
						end

						10'h10: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp51) ? 10'h14 : 10'h44);

									end
								end

							endcase
						end

						10'h11: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h10;

									end
								end

							endcase
						end

						10'h14: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h15;

									end
								end

							endcase
						end

						10'h15: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp55) ? 10'h18 : 10'h1a);

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h15;

									end
								end

							endcase
						end

						10'h1a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1b;

									end
								end

							endcase
						end

						10'h1b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp130) ? 10'h1e : 10'h20);

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1b;

									end
								end

							endcase
						end

						10'h20: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h21;

									end
								end

							endcase
						end

						10'h21: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp219) ? 10'h24 : 10'h26);

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h21;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h27;

									end
								end

							endcase
						end

						10'h27: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp308) ? 10'h2a : 10'h2c);

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h27;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h2d;

									end
								end

							endcase
						end

						10'h2d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp397) ? 10'h30 : 10'h32);

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h2d;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h33;

									end
								end

							endcase
						end

						10'h33: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp486) ? 10'h36 : 10'h38);

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h33;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h39;

									end
								end

							endcase
						end

						10'h39: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp575) ? 10'h3c : 10'h3e);

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h39;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h3f;

									end
								end

							endcase
						end

						10'h3f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp664) ? 10'h42 : 10'h11);

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h3f;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h45;

									end
								end

							endcase
						end

						10'h45: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp753) ? 10'h49 : 10'h79);

									end
								end

							endcase
						end

						10'h46: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h45;

									end
								end

							endcase
						end

						10'h49: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h4a;

									end
								end

							endcase
						end

						10'h4a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp757) ? 10'h4d : 10'h4f);

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h4a;

									end
								end

							endcase
						end

						10'h4f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h50;

									end
								end

							endcase
						end

						10'h50: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp832) ? 10'h53 : 10'h55);

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h50;

									end
								end

							endcase
						end

						10'h55: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h56;

									end
								end

							endcase
						end

						10'h56: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp921) ? 10'h59 : 10'h5b);

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h56;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h5c;

									end
								end

							endcase
						end

						10'h5c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1010) ? 10'h5f : 10'h61);

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h5c;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h62;

									end
								end

							endcase
						end

						10'h62: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1099) ? 10'h65 : 10'h67);

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h62;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h68;

									end
								end

							endcase
						end

						10'h68: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1188) ? 10'h6b : 10'h6d);

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h68;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h6e;

									end
								end

							endcase
						end

						10'h6e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1277) ? 10'h71 : 10'h73);

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h6e;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h74;

									end
								end

							endcase
						end

						10'h74: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1366) ? 10'h77 : 10'h46);

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h74;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h7a;

									end
								end

							endcase
						end

						10'h7a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1455) ? 10'h7e : 10'hae);

									end
								end

							endcase
						end

						10'h7b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h7a;

									end
								end

							endcase
						end

						10'h7e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h7f;

									end
								end

							endcase
						end

						10'h7f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1459) ? 10'h82 : 10'h84);

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h7f;

									end
								end

							endcase
						end

						10'h84: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h85;

									end
								end

							endcase
						end

						10'h85: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1534) ? 10'h88 : 10'h8a);

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h85;

									end
								end

							endcase
						end

						10'h8a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h8b;

									end
								end

							endcase
						end

						10'h8b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1623) ? 10'h8e : 10'h90);

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h8b;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h91;

									end
								end

							endcase
						end

						10'h91: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1712) ? 10'h94 : 10'h96);

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h91;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h97;

									end
								end

							endcase
						end

						10'h97: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1801) ? 10'h9a : 10'h9c);

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h97;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h9d;

									end
								end

							endcase
						end

						10'h9d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1890) ? 10'ha0 : 10'ha2);

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h9d;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'ha3;

									end
								end

							endcase
						end

						10'ha3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1979) ? 10'ha6 : 10'ha8);

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'ha3;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'ha9;

									end
								end

							endcase
						end

						10'ha9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2068) ? 10'hac : 10'h7b);

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'ha9;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'haf;

									end
								end

							endcase
						end

						10'haf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2157) ? 10'hb3 : 10'he3);

									end
								end

							endcase
						end

						10'hb0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'haf;

									end
								end

							endcase
						end

						10'hb3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hb4;

									end
								end

							endcase
						end

						10'hb4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2161) ? 10'hb7 : 10'hb9);

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hb4;

									end
								end

							endcase
						end

						10'hb9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hba;

									end
								end

							endcase
						end

						10'hba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2236) ? 10'hbd : 10'hbf);

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hba;

									end
								end

							endcase
						end

						10'hbf: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hc0;

									end
								end

							endcase
						end

						10'hc0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2325) ? 10'hc3 : 10'hc5);

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hc0;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hc6;

									end
								end

							endcase
						end

						10'hc6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2414) ? 10'hc9 : 10'hcb);

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hc6;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hcc;

									end
								end

							endcase
						end

						10'hcc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2503) ? 10'hcf : 10'hd1);

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hcc;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hd2;

									end
								end

							endcase
						end

						10'hd2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2592) ? 10'hd5 : 10'hd7);

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hd2;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hd8;

									end
								end

							endcase
						end

						10'hd8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2681) ? 10'hdb : 10'hdd);

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hd8;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hde;

									end
								end

							endcase
						end

						10'hde: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2770) ? 10'he1 : 10'hb0);

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'hde;

									end
								end

							endcase
						end

						10'he3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'he4;

									end
								end

							endcase
						end

						10'he4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2858) ? 10'he7 : 10'h133);

									end
								end

							endcase
						end

						10'he5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'he4;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h1e: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 10'he9;

									end
								end

							endcase
						end

						10'he9: begin

							case(r_sys_run_stage) 
								6'h1f: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_phase <= 10'heb;

									end
								end

							endcase
						end

						10'heb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hec;

									end
								end

							endcase
						end

						10'hec: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2862) ? 10'hef : 10'hf1);

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'hec;

									end
								end

							endcase
						end

						10'hf1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hf2;

									end
								end

							endcase
						end

						10'hf2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2946) ? 10'hf5 : 10'hf7);

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'hf2;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hf8;

									end
								end

							endcase
						end

						10'hf8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3030) ? 10'hfb : 10'hfd);

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'hf8;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'hfe;

									end
								end

							endcase
						end

						10'hfe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3114) ? 10'h101 : 10'h103);

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_phase <= 10'hfe;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h104;

									end
								end

							endcase
						end

						10'h104: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3197) ? 10'h107 : 10'h109);

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h104;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h10a;

									end
								end

							endcase
						end

						10'h10a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp3698) ? 10'h10d : 10'h10f);

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h10a;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h110;

									end
								end

							endcase
						end

						10'h110: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4199) ? 10'h113 : 10'h115);

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h110;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h116;

									end
								end

							endcase
						end

						10'h116: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp4700) ? 10'h119 : 10'h11b);

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h116;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h11c;

									end
								end

							endcase
						end

						10'h11c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5201) ? 10'h11f : 10'h121);

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h11c;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h122;

									end
								end

							endcase
						end

						10'h122: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5702) ? 10'h125 : 10'h127);

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h122;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h128;

									end
								end

							endcase
						end

						10'h128: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6203) ? 10'h12b : 10'h12d);

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_phase <= 10'h128;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h12e;

									end
								end

							endcase
						end

						10'h12e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp6704) ? 10'h131 : 10'he5);

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3a)) begin
										r_sys_run_phase <= 10'h12e;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h134;

									end
								end

							endcase
						end

						10'h134: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7193) ? 10'h138 : 10'h168);

									end
								end

							endcase
						end

						10'h135: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h134;

									end
								end

							endcase
						end

						10'h138: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h139;

									end
								end

							endcase
						end

						10'h139: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7198) ? 10'h13c : 10'h13e);

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h139;

									end
								end

							endcase
						end

						10'h13e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h13f;

									end
								end

							endcase
						end

						10'h13f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7273) ? 10'h142 : 10'h144);

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h13f;

									end
								end

							endcase
						end

						10'h144: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h145;

									end
								end

							endcase
						end

						10'h145: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7369) ? 10'h148 : 10'h14a);

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h145;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h14b;

									end
								end

							endcase
						end

						10'h14b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7465) ? 10'h14e : 10'h150);

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h14b;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h151;

									end
								end

							endcase
						end

						10'h151: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7561) ? 10'h154 : 10'h156);

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h151;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h157;

									end
								end

							endcase
						end

						10'h157: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7657) ? 10'h15a : 10'h15c);

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h157;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h15d;

									end
								end

							endcase
						end

						10'h15d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7753) ? 10'h160 : 10'h162);

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h15d;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h163;

									end
								end

							endcase
						end

						10'h163: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7849) ? 10'h166 : 10'h135);

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h163;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h169;

									end
								end

							endcase
						end

						10'h169: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7945) ? 10'h16d : 10'h19d);

									end
								end

							endcase
						end

						10'h16a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h169;

									end
								end

							endcase
						end

						10'h16d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h16e;

									end
								end

							endcase
						end

						10'h16e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7950) ? 10'h171 : 10'h173);

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h16e;

									end
								end

							endcase
						end

						10'h173: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h174;

									end
								end

							endcase
						end

						10'h174: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8025) ? 10'h177 : 10'h179);

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h174;

									end
								end

							endcase
						end

						10'h179: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h17a;

									end
								end

							endcase
						end

						10'h17a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8121) ? 10'h17d : 10'h17f);

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h17a;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h180;

									end
								end

							endcase
						end

						10'h180: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8217) ? 10'h183 : 10'h185);

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h180;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h186;

									end
								end

							endcase
						end

						10'h186: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8313) ? 10'h189 : 10'h18b);

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h186;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h18c;

									end
								end

							endcase
						end

						10'h18c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8409) ? 10'h18f : 10'h191);

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h18c;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h192;

									end
								end

							endcase
						end

						10'h192: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8505) ? 10'h195 : 10'h197);

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h192;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h198;

									end
								end

							endcase
						end

						10'h198: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8601) ? 10'h19b : 10'h16a);

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h198;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h19e;

									end
								end

							endcase
						end

						10'h19e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8697) ? 10'h1a2 : 10'h1d2);

									end
								end

							endcase
						end

						10'h19f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h19e;

									end
								end

							endcase
						end

						10'h1a2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1a3;

									end
								end

							endcase
						end

						10'h1a3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8702) ? 10'h1a6 : 10'h1a8);

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1a3;

									end
								end

							endcase
						end

						10'h1a8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1a9;

									end
								end

							endcase
						end

						10'h1a9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8777) ? 10'h1ac : 10'h1ae);

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1a9;

									end
								end

							endcase
						end

						10'h1ae: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1af;

									end
								end

							endcase
						end

						10'h1af: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8873) ? 10'h1b2 : 10'h1b4);

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1af;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1b5;

									end
								end

							endcase
						end

						10'h1b5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp8969) ? 10'h1b8 : 10'h1ba);

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1b5;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1bb;

									end
								end

							endcase
						end

						10'h1bb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9065) ? 10'h1be : 10'h1c0);

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1bb;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1c1;

									end
								end

							endcase
						end

						10'h1c1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9161) ? 10'h1c4 : 10'h1c6);

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1c1;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1c7;

									end
								end

							endcase
						end

						10'h1c7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9257) ? 10'h1ca : 10'h1cc);

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1c7;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1cd;

									end
								end

							endcase
						end

						10'h1cd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9353) ? 10'h1d0 : 10'h19f);

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1cd;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1d3;

									end
								end

							endcase
						end

						10'h1d3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9449) ? 10'h1d7 : 10'h207);

									end
								end

							endcase
						end

						10'h1d4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1d3;

									end
								end

							endcase
						end

						10'h1d7: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1d8;

									end
								end

							endcase
						end

						10'h1d8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9454) ? 10'h1db : 10'h1dd);

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1d8;

									end
								end

							endcase
						end

						10'h1dd: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1de;

									end
								end

							endcase
						end

						10'h1de: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9529) ? 10'h1e1 : 10'h1e3);

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1de;

									end
								end

							endcase
						end

						10'h1e3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1e4;

									end
								end

							endcase
						end

						10'h1e4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9625) ? 10'h1e7 : 10'h1e9);

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1e4;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1ea;

									end
								end

							endcase
						end

						10'h1ea: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9721) ? 10'h1ed : 10'h1ef);

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1ea;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1f0;

									end
								end

							endcase
						end

						10'h1f0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9817) ? 10'h1f3 : 10'h1f5);

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1f0;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1f6;

									end
								end

							endcase
						end

						10'h1f6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp9913) ? 10'h1f9 : 10'h1fb);

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1f6;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h1fc;

									end
								end

							endcase
						end

						10'h1fc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10009) ? 10'h1ff : 10'h201);

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h1fc;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= 10'h202;

									end
								end

							endcase
						end

						10'h202: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10105) ? 10'h205 : 10'h1d4);

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_phase <= 10'h202;

									end
								end

							endcase
						end

						10'h207: begin
							r_sys_run_phase <= 10'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h10: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h11: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h14: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h15: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h20: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h21: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h27: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h2d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h33: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h39: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h3f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h45: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h46: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h49: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h4a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h4f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h50: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h55: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h56: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h5c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h62: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h68: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h6e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h74: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h7a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h7b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h7e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h7f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h84: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h85: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h8a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h8b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h91: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h97: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h9d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'ha9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'haf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hb0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hb3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hb4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hb9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hbf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hcc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hd8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hde: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'he9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1f: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'heb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hec: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hf8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'hfe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h104: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h10a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h110: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h116: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h11c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h122: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h128: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h12e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3a)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h134: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h135: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h138: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h139: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h13e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h13f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h144: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h145: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h14b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h151: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h157: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h15d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h163: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h169: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h16a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h16d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h16e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h173: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h174: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h179: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h17a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h180: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h186: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h18c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h192: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h198: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h19e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h19f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1a9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ae: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1af: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1bb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1c7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1cd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1d8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1dd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1de: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ea: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1fc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h202: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_stage <= 6'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 6'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h11: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h14: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h20: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h21: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h27: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h2d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h33: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h39: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h3f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h45: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h46: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h49: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h4a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h4f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h50: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h55: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h56: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h62: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h68: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h6e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h74: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h7a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h7b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h7e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h7f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h84: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h85: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h8a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h8b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h91: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h97: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h9d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'ha9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'haf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hb9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hbf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hcc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hd8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hde: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'he9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub16_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub17_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub18_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub19_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub20_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub21_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub22_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub23_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub24_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub25_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub26_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub27_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub28_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub29_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub30_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1f: begin
									if((r_sys_run_step==6'h1)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= ((w_sub31_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						10'heb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hec: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hf8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'hfe: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h1c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h104: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h110: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h116: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h11c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h122: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h128: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h3c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h3d)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h12e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3a)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h39)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h134: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h135: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h138: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h139: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h13e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h13f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h144: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h145: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h14b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h151: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h157: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h15d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h163: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h169: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h16a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h16d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h16e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h173: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h174: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h179: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h17a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h180: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h186: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h18c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h192: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h198: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h19e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h19f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1a9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1ae: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1af: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1bb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1c7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1cd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1d8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1dd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1de: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1e3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ea: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1fc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
									else
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h202: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==6'h8)) begin
										r_sys_run_step <= 6'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						10'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						10'h207: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_addr_1 <= 15'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp10[14:0] );

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp64[14:0] );

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp141[14:0] );

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp230[14:0] );

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp319[14:0] );

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp408[14:0] );

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp497[14:0] );

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp586[14:0] );

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp675[14:0] );

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp766[14:0] );

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp843[14:0] );

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp932[14:0] );

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1021[14:0] );

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1110[14:0] );

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1199[14:0] );

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1288[14:0] );

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1377[14:0] );

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1468[14:0] );

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1545[14:0] );

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1634[14:0] );

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1723[14:0] );

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1812[14:0] );

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1901[14:0] );

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp1990[14:0] );

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2079[14:0] );

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2170[14:0] );

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2247[14:0] );

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2336[14:0] );

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2425[14:0] );

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2514[14:0] );

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2603[14:0] );

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2692[14:0] );

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp2781[14:0] );

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp7203[14:0] );

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp7280[14:0] );

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp7376[14:0] );

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp7472[14:0] );

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp7568[14:0] );

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp7664[14:0] );

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp7760[14:0] );

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp7856[14:0] );

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp7955[14:0] );

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8032[14:0] );

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8128[14:0] );

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8224[14:0] );

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8320[14:0] );

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8416[14:0] );

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8512[14:0] );

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8608[14:0] );

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8707[14:0] );

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8784[14:0] );

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8880[14:0] );

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp8976[14:0] );

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp9072[14:0] );

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp9168[14:0] );

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp9264[14:0] );

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp9360[14:0] );

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp9459[14:0] );

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp9536[14:0] );

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp9632[14:0] );

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp9728[14:0] );

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp9824[14:0] );

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp9920[14:0] );

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp10016[14:0] );

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_addr_1 <= $signed( w_sys_tmp10112[14:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp13;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp7206;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp7283;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp7379;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp7475;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp7571;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp7667;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp7763;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp7859;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp7958;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8035;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8131;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8227;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8323;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8419;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8515;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8611;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8710;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8787;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8883;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp8979;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp9075;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp9171;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp9267;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp9363;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp9462;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp9539;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp9635;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp9731;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp9827;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp9923;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp10019;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_datain_1 <= w_sys_tmp10115;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_u_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_fld_u_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h207: begin
							r_fld_u_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp5;

									end
								end

							endcase
						end

						10'hf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h11: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp54;

									end
								end

							endcase
						end

						10'h44: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp752;

									end
								end

							endcase
						end

						10'h46: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp756;

									end
								end

							endcase
						end

						10'h79: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp1454;

									end
								end

							endcase
						end

						10'h7b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp1458;

									end
								end

							endcase
						end

						10'hae: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp2156;

									end
								end

							endcase
						end

						10'hb0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp2160;

									end
								end

							endcase
						end

						10'heb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp2861;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_33 <= w_sys_tmp2944;

									end
								end

							endcase
						end

						10'hf1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp2945;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_33 <= w_sys_tmp3028;

									end
								end

							endcase
						end

						10'hf7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp3029;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_33 <= w_sys_tmp3112;

									end
								end

							endcase
						end

						10'hfd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp3113;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_run_k_33 <= w_sys_tmp3196;

									end
								end

							endcase
						end

						10'h133: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp7192;

									end
								end

							endcase
						end

						10'h135: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp7196;

									end
								end

							endcase
						end

						10'h168: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp7944;

									end
								end

							endcase
						end

						10'h16a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp7948;

									end
								end

							endcase
						end

						10'h19d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp8696;

									end
								end

							endcase
						end

						10'h19f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp8700;

									end
								end

							endcase
						end

						10'h1d2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp9448;

									end
								end

							endcase
						end

						10'h1d4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_k_33 <= w_sys_tmp9452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'hd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp14;

									end
								end

							endcase
						end

						10'h14: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_34 <= w_sys_tmp68;

									end
								end

							endcase
						end

						10'h1a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp129;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp145;

									end
								end

							endcase
						end

						10'h20: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp218;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp234;

									end
								end

							endcase
						end

						10'h26: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp307;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp323;

									end
								end

							endcase
						end

						10'h2c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp396;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp412;

									end
								end

							endcase
						end

						10'h32: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp485;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp501;

									end
								end

							endcase
						end

						10'h38: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp574;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp590;

									end
								end

							endcase
						end

						10'h3e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp663;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp679;

									end
								end

							endcase
						end

						10'h49: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_34 <= w_sys_tmp770;

									end
								end

							endcase
						end

						10'h4f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp831;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp847;

									end
								end

							endcase
						end

						10'h55: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp920;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp936;

									end
								end

							endcase
						end

						10'h5b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1009;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1025;

									end
								end

							endcase
						end

						10'h61: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1098;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1114;

									end
								end

							endcase
						end

						10'h67: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1187;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1203;

									end
								end

							endcase
						end

						10'h6d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1276;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1292;

									end
								end

							endcase
						end

						10'h73: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1365;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1381;

									end
								end

							endcase
						end

						10'h7e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_34 <= w_sys_tmp1472;

									end
								end

							endcase
						end

						10'h84: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1533;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1549;

									end
								end

							endcase
						end

						10'h8a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1622;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1638;

									end
								end

							endcase
						end

						10'h90: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1711;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1727;

									end
								end

							endcase
						end

						10'h96: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1800;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1816;

									end
								end

							endcase
						end

						10'h9c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1889;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1905;

									end
								end

							endcase
						end

						10'ha2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp1978;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp1994;

									end
								end

							endcase
						end

						10'ha8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp2067;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp2083;

									end
								end

							endcase
						end

						10'hb3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_34 <= w_sys_tmp2174;

									end
								end

							endcase
						end

						10'hb9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp2235;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp2251;

									end
								end

							endcase
						end

						10'hbf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp2324;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp2340;

									end
								end

							endcase
						end

						10'hc5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp2413;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp2429;

									end
								end

							endcase
						end

						10'hcb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp2502;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp2518;

									end
								end

							endcase
						end

						10'hd1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp2591;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp2607;

									end
								end

							endcase
						end

						10'hd7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp2680;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp2696;

									end
								end

							endcase
						end

						10'hdd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp2769;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_j_34 <= w_sys_tmp2785;

									end
								end

							endcase
						end

						10'h103: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_34 <= w_sys_tmp3270;

									end
								end

							endcase
						end

						10'h109: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp3697;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_34 <= w_sys_tmp3771;

									end
								end

							endcase
						end

						10'h10f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp4198;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_34 <= w_sys_tmp4272;

									end
								end

							endcase
						end

						10'h115: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp4699;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_34 <= w_sys_tmp4773;

									end
								end

							endcase
						end

						10'h11b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp5200;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_34 <= w_sys_tmp5274;

									end
								end

							endcase
						end

						10'h121: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp5701;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_34 <= w_sys_tmp5775;

									end
								end

							endcase
						end

						10'h127: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp6202;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_34 <= w_sys_tmp6276;

									end
								end

							endcase
						end

						10'h12d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp6703;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_run_j_34 <= w_sys_tmp6777;

									end
								end

							endcase
						end

						10'h138: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp7197;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_34 <= w_sys_tmp7211;

									end
								end

							endcase
						end

						10'h13e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp7272;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp7289;

									end
								end

							endcase
						end

						10'h144: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp7368;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp7385;

									end
								end

							endcase
						end

						10'h14a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp7464;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp7481;

									end
								end

							endcase
						end

						10'h150: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp7560;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp7577;

									end
								end

							endcase
						end

						10'h156: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp7656;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp7673;

									end
								end

							endcase
						end

						10'h15c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp7752;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp7769;

									end
								end

							endcase
						end

						10'h162: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp7848;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp7865;

									end
								end

							endcase
						end

						10'h16d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp7949;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_34 <= w_sys_tmp7963;

									end
								end

							endcase
						end

						10'h173: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8024;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp8041;

									end
								end

							endcase
						end

						10'h179: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8120;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp8137;

									end
								end

							endcase
						end

						10'h17f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8216;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp8233;

									end
								end

							endcase
						end

						10'h185: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8312;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp8329;

									end
								end

							endcase
						end

						10'h18b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8408;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp8425;

									end
								end

							endcase
						end

						10'h191: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8504;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp8521;

									end
								end

							endcase
						end

						10'h197: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8600;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp8617;

									end
								end

							endcase
						end

						10'h1a2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8701;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_34 <= w_sys_tmp8715;

									end
								end

							endcase
						end

						10'h1a8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8776;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp8793;

									end
								end

							endcase
						end

						10'h1ae: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8872;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp8889;

									end
								end

							endcase
						end

						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp8968;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp8985;

									end
								end

							endcase
						end

						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp9064;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp9081;

									end
								end

							endcase
						end

						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp9160;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp9177;

									end
								end

							endcase
						end

						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp9256;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp9273;

									end
								end

							endcase
						end

						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp9352;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp9369;

									end
								end

							endcase
						end

						10'h1d7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp9453;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_j_34 <= w_sys_tmp9467;

									end
								end

							endcase
						end

						10'h1dd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp9528;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp9545;

									end
								end

							endcase
						end

						10'h1e3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp9624;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp9641;

									end
								end

							endcase
						end

						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp9720;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp9737;

									end
								end

							endcase
						end

						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp9816;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp9833;

									end
								end

							endcase
						end

						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp9912;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp9929;

									end
								end

							endcase
						end

						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp10008;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp10025;

									end
								end

							endcase
						end

						10'h201: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_j_34 <= w_sys_tmp10104;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_j_34 <= w_sys_tmp10121;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_35 <= w_sys_intOne;

									end
								end

							endcase
						end

						10'he5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_n_35 <= w_sys_tmp2860;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_mx_36 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_my_37 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_nlast_38 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp134;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp223;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp312;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp401;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp490;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp579;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp668;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp836;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp925;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1014;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1103;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1192;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1281;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1370;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1538;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1627;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1716;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1805;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1894;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp1983;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp2072;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp2240;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp2329;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp2418;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp2507;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp2596;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp2685;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (6'h2<=r_sys_run_step && r_sys_run_step<=6'h7)) begin
										r_run_tmpj_39 <= w_sys_tmp2774;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp7277;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp7373;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp7469;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp7565;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp7661;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp7757;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp7853;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp8029;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp8125;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp8221;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp8317;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp8413;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp8509;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp8605;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp8781;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp8877;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp8973;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp9069;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp9165;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp9261;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp9357;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp9533;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp9629;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp9725;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp9821;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp9917;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp10013;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_tmpj_39 <= w_sys_tmp10109;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_40 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h18: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_40 <= w_sys_tmp67;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_41 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_41 <= w_sys_tmp144;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h20: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_42 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_42 <= w_sys_tmp233;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h26: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_43 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_43 <= w_sys_tmp322;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_44 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_44 <= w_sys_tmp411;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h32: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_45 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_45 <= w_sys_tmp500;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h38: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_46 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_46 <= w_sys_tmp589;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_47 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_47 <= w_sys_tmp678;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h49: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_48 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h4d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_48 <= w_sys_tmp769;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_49 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_49 <= w_sys_tmp846;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h55: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_50 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_50 <= w_sys_tmp935;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_51 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_51 <= w_sys_tmp1024;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h61: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_52 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_52 <= w_sys_tmp1113;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h67: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_53 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_53 <= w_sys_tmp1202;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_54 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_54 <= w_sys_tmp1291;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h73: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_55 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_55 <= w_sys_tmp1380;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h7e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_56 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h82: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_56 <= w_sys_tmp1471;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h84: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_57 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_57 <= w_sys_tmp1548;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_58 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_58 <= w_sys_tmp1637;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h90: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_59 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_59 <= w_sys_tmp1726;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h96: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_60 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_60 <= w_sys_tmp1815;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_61 <= r_run_j_34;

									end
								end

							endcase
						end

						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_61 <= w_sys_tmp1904;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_62 <= r_run_j_34;

									end
								end

							endcase
						end

						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_62 <= w_sys_tmp1993;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_63 <= r_run_j_34;

									end
								end

							endcase
						end

						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_63 <= w_sys_tmp2082;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_64 <= r_run_j_34;

									end
								end

							endcase
						end

						10'hb7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_64 <= w_sys_tmp2173;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_65 <= r_run_j_34;

									end
								end

							endcase
						end

						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_65 <= w_sys_tmp2250;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbf: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_66 <= r_run_j_34;

									end
								end

							endcase
						end

						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_66 <= w_sys_tmp2339;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_67 <= r_run_j_34;

									end
								end

							endcase
						end

						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_67 <= w_sys_tmp2428;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_68 <= r_run_j_34;

									end
								end

							endcase
						end

						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_68 <= w_sys_tmp2517;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd1: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_69 <= r_run_j_34;

									end
								end

							endcase
						end

						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_69 <= w_sys_tmp2606;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd7: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_70 <= r_run_j_34;

									end
								end

							endcase
						end

						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_70 <= w_sys_tmp2695;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdd: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_71 <= r_run_j_34;

									end
								end

							endcase
						end

						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_71 <= w_sys_tmp2784;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_72 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_72 <= w_sys_tmp3259;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_73 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_73 <= w_sys_tmp3260;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_74 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_74 <= w_sys_tmp3261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_75 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_75 <= w_sys_tmp3262;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_76 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_76 <= w_sys_tmp3263;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_77 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_77 <= w_sys_tmp3264;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_78 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_78 <= w_sys_tmp3265;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_79 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_79 <= w_sys_tmp3266;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_80 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_80 <= w_sys_tmp3267;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_81 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_81 <= w_sys_tmp3268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h103: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_82 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_82 <= w_sys_tmp3269;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_83 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_83 <= w_sys_tmp3760;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_84 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_84 <= w_sys_tmp3761;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_85 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_85 <= w_sys_tmp3762;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_86 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_86 <= w_sys_tmp3763;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_87 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_87 <= w_sys_tmp3764;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_88 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_88 <= w_sys_tmp3765;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_89 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_89 <= w_sys_tmp3766;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_90 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_90 <= w_sys_tmp3767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_91 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_91 <= w_sys_tmp3768;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_92 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_92 <= w_sys_tmp3769;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h109: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_93 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_93 <= w_sys_tmp3770;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_94 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_94 <= w_sys_tmp4261;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_95 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_95 <= w_sys_tmp4262;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_96 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_96 <= w_sys_tmp4263;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_97 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_97 <= w_sys_tmp4264;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_98 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_98 <= w_sys_tmp4265;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_99 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_99 <= w_sys_tmp4266;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_100 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_100 <= w_sys_tmp4267;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_101 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_101 <= w_sys_tmp4268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_102 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_102 <= w_sys_tmp4269;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_103 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_103 <= w_sys_tmp4270;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h10f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_104 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_104 <= w_sys_tmp4271;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_105 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_105 <= w_sys_tmp4762;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_106 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_106 <= w_sys_tmp4763;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_107 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_107 <= w_sys_tmp4764;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_108 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_108 <= w_sys_tmp4765;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_109 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_109 <= w_sys_tmp4766;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_110 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_110 <= w_sys_tmp4767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_111 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_111 <= w_sys_tmp4768;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_112 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_112 <= w_sys_tmp4769;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_113 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_113 <= w_sys_tmp4770;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_114 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_114 <= w_sys_tmp4771;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h115: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_115 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_115 <= w_sys_tmp4772;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_116 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_116 <= w_sys_tmp5263;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_117 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_117 <= w_sys_tmp5264;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_118 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_118 <= w_sys_tmp5265;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_119 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_119 <= w_sys_tmp5266;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_120 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_120 <= w_sys_tmp5267;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_121 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_121 <= w_sys_tmp5268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_122 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_122 <= w_sys_tmp5269;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_123 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_123 <= w_sys_tmp5270;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_124 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_124 <= w_sys_tmp5271;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_125 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_125 <= w_sys_tmp5272;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h11b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_126 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_126 <= w_sys_tmp5273;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_127 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_127 <= w_sys_tmp5764;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_128 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_128 <= w_sys_tmp5765;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_129 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_129 <= w_sys_tmp5766;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_130 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_130 <= w_sys_tmp5767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_131 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_131 <= w_sys_tmp5768;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_132 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_132 <= w_sys_tmp5769;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_133 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_133 <= w_sys_tmp5770;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_134 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_134 <= w_sys_tmp5771;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_135 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_135 <= w_sys_tmp5772;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_136 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_136 <= w_sys_tmp5773;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h121: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_137 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_137 <= w_sys_tmp5774;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_138 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_run_copy0_j_138 <= w_sys_tmp6265;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_139 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_run_copy1_j_139 <= w_sys_tmp6266;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_140 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy2_j_140 <= w_sys_tmp6267;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_141 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_141 <= w_sys_tmp6268;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_142 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_142 <= w_sys_tmp6269;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_143 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_143 <= w_sys_tmp6270;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_144 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_run_copy6_j_144 <= w_sys_tmp6271;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_145 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_145 <= w_sys_tmp6272;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_146 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_146 <= w_sys_tmp6273;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_147 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_147 <= w_sys_tmp6274;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h127: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_148 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_148 <= w_sys_tmp6275;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_149 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_149 <= w_sys_tmp6766;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_150 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'he)) begin
										r_run_copy1_j_150 <= w_sys_tmp6767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy2_j_151 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_run_copy2_j_151 <= w_sys_tmp6768;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy3_j_152 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_run_copy3_j_152 <= w_sys_tmp6769;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy4_j_153 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_run_copy4_j_153 <= w_sys_tmp6770;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy5_j_154 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_run_copy5_j_154 <= w_sys_tmp6771;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy6_j_155 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy6_j_155 <= w_sys_tmp6772;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy7_j_156 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_run_copy7_j_156 <= w_sys_tmp6773;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy8_j_157 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_run_copy8_j_157 <= w_sys_tmp6774;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy9_j_158 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_run_copy9_j_158 <= w_sys_tmp6775;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h12d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy10_j_159 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_run_copy10_j_159 <= w_sys_tmp6776;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h138: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_160 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_160 <= w_sys_tmp7210;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_161 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_161 <= w_sys_tmp7287;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h13e: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_162 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_162 <= w_sys_tmp7288;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h144: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_163 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_163 <= w_sys_tmp7383;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h144: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_164 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_164 <= w_sys_tmp7384;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_165 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_165 <= w_sys_tmp7479;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h14a: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_166 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_166 <= w_sys_tmp7480;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h150: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_167 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_167 <= w_sys_tmp7575;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h150: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_168 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_168 <= w_sys_tmp7576;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h156: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_169 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_169 <= w_sys_tmp7671;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h156: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_170 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_170 <= w_sys_tmp7672;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h15c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_171 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_171 <= w_sys_tmp7767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h15c: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_172 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_172 <= w_sys_tmp7768;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h162: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_173 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_173 <= w_sys_tmp7863;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h162: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_174 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_174 <= w_sys_tmp7864;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h16d: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_175 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_175 <= w_sys_tmp7962;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h173: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_176 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_176 <= w_sys_tmp8039;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h173: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_177 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_177 <= w_sys_tmp8040;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h179: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_178 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_178 <= w_sys_tmp8135;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h179: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_179 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_179 <= w_sys_tmp8136;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h17f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_180 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_180 <= w_sys_tmp8231;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h17f: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_181 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_181 <= w_sys_tmp8232;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h185: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_182 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_182 <= w_sys_tmp8327;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h185: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_183 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_183 <= w_sys_tmp8328;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_184 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_184 <= w_sys_tmp8423;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18b: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_185 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_185 <= w_sys_tmp8424;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h191: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_186 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_186 <= w_sys_tmp8519;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h191: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_187 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_187 <= w_sys_tmp8520;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h197: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_188 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_188 <= w_sys_tmp8615;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h197: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_189 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_189 <= w_sys_tmp8616;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a2: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_190 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_190 <= w_sys_tmp8714;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_191 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_191 <= w_sys_tmp8791;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1a8: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_192 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_192 <= w_sys_tmp8792;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ae: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_193 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_193 <= w_sys_tmp8887;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ae: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_194 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_194 <= w_sys_tmp8888;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_195 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_195 <= w_sys_tmp8983;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1b4: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_196 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_196 <= w_sys_tmp8984;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_197 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_197 <= w_sys_tmp9079;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ba: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_198 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_198 <= w_sys_tmp9080;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_199 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_199 <= w_sys_tmp9175;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c0: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_200 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_200 <= w_sys_tmp9176;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_201 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_201 <= w_sys_tmp9271;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1c6: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_202 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_202 <= w_sys_tmp9272;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_203 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_203 <= w_sys_tmp9367;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1cc: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_204 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_204 <= w_sys_tmp9368;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1d7: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_205 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_205 <= w_sys_tmp9466;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1dd: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_206 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_206 <= w_sys_tmp9543;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1dd: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_207 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_207 <= w_sys_tmp9544;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_208 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_208 <= w_sys_tmp9639;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e3: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_209 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_209 <= w_sys_tmp9640;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_210 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_210 <= w_sys_tmp9735;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e9: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_211 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_211 <= w_sys_tmp9736;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_212 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_212 <= w_sys_tmp9831;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1ef: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_213 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_213 <= w_sys_tmp9832;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_214 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_214 <= w_sys_tmp9927;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1f5: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_215 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_215 <= w_sys_tmp9928;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_216 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_216 <= w_sys_tmp10023;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1fb: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_217 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_217 <= w_sys_tmp10024;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h201: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy0_j_218 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_run_copy0_j_218 <= w_sys_tmp10119;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h201: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_run_copy1_j_219 <= r_run_j_34;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_run_copy1_j_219 <= w_sys_tmp10120;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h12: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_u_addr <= $signed( w_sys_tmp1719[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_u_datain <= w_sys_tmp1722;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h94: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub19_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub19_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp3047[11:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp3035[11:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp3041[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp3038[11:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4744[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4734[11:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4758[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp4729[11:0] );

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp8980[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub19_result_datain <= w_sys_tmp3065;

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub19_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub19_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub19_result_datain <= w_sys_tmp4709;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1) || (r_sys_run_step==6'hf)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub19_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub19_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1b8: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub19_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'hb: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_u_addr <= $signed( w_sys_tmp1106[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_u_datain <= w_sys_tmp1109;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h65: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub12_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub12_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp2963[11:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp2951[11:0] );

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp2957[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp2954[11:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5211[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5226[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5240[11:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp5216[11:0] );

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp8324[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_sub12_result_datain <= w_sys_tmp2992;

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub12_result_datain <= r_sys_tmp2_float;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub12_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub12_result_datain <= w_sys_tmp5258;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub12_result_datain <= w_sys_tmp5220;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub12_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h189: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'ha: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_u_addr <= $signed( w_sys_tmp1017[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_u_datain <= w_sys_tmp1020;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h5f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub11_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub11_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp2963[11:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp2951[11:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp2957[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp2954[11:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4739[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4725[11:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4715[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp4710[11:0] );

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp8228[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub11_result_datain <= w_sys_tmp2981;

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub11_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub11_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_datain <= w_sys_tmp4757;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub11_result_datain <= w_sys_tmp4719;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hf)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub11_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h183: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'hd: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_u_addr <= $signed( w_sys_tmp1284[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_u_datain <= w_sys_tmp1287;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h71: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub14_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub14_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2963[11:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2951[11:0] );

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2957[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp2954[11:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp6218[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp6242[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp6213[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp6228[11:0] );

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp8516[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub14_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub14_result_datain <= w_sys_tmp3014;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub14_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub14_result_datain <= w_sys_tmp6260;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub14_result_datain <= w_sys_tmp6222;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub14_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h195: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'hc: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_u_addr <= $signed( w_sys_tmp1195[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_u_datain <= w_sys_tmp1198;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h6b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub13_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub13_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2963[11:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2951[11:0] );

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2957[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp2954[11:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5717[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5741[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5727[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp5712[11:0] );

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp8420[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub13_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub13_result_datain <= w_sys_tmp3003;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_datain <= w_sys_tmp5759;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub13_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub13_result_datain <= w_sys_tmp5721;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub13_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h18f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'hf: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_u_addr <= $signed( w_sys_tmp1464[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_u_datain <= w_sys_tmp1467;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h82: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub16_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub16_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp3044[11:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp3035[11:0] );

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp3226[11:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp3255[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp3241[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp3231[11:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp6762[11:0] );

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp8711[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub16_result_datain <= w_sys_tmp3037;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub16_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub16_result_datain <= w_sys_tmp3206;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub16_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub16_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h1a6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub16_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'he: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_u_addr <= $signed( w_sys_tmp1373[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_u_datain <= w_sys_tmp1376;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h77: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub15_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub15_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp2957[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp2954[11:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6714[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6743[11:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6719[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp6729[11:0] );

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp8612[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub15_result_datain <= w_sys_tmp3025;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub15_result_datain <= w_sys_tmp6723;

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_datain <= r_sys_tmp7_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub15_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h19b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h11: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_u_addr <= $signed( w_sys_tmp1630[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_u_datain <= w_sys_tmp1633;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h8e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub18_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub18_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp3047[11:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp3035[11:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp3041[11:0] );

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4228[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4233[11:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4257[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp4243[11:0] );

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp8884[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub18_result_datain <= w_sys_tmp3037;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub18_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub18_result_datain <= w_sys_tmp4208;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub18_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub18_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub18_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1b2: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub18_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h10: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_u_addr <= $signed( w_sys_tmp1541[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_u_datain <= w_sys_tmp1544;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h88: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub17_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub17_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3047[11:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3035[11:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3041[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3038[11:0] );

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3756[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3727[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3742[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp3732[11:0] );

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp8788[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub17_result_datain <= w_sys_tmp3043;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub17_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub17_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub17_result_datain <= w_sys_tmp3707;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub17_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub17_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub17_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h13: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub20_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub20_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_u_addr <= $signed( w_sys_tmp1808[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_u_datain <= w_sys_tmp1811;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h9a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub20_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub20_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp3047[11:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp3035[11:0] );

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp3041[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp3038[11:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp5259[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp5235[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp5245[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp5230[11:0] );

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp9076[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_sub20_result_datain <= w_sys_tmp3076;

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub20_result_datain <= r_sys_tmp2_float;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub20_result_datain <= w_sys_tmp5210;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub20_result_datain <= r_sys_tmp0_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub20_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub20_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1be: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub20_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h14: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub21_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub21_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_u_addr <= $signed( w_sys_tmp1897[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_u_datain <= w_sys_tmp1900;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub21_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub21_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp3047[11:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp3035[11:0] );

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp3041[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp3038[11:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp5731[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp5746[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp5736[11:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp5760[11:0] );

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp9172[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub21_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub21_result_datain <= w_sys_tmp3087;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub21_result_datain <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub21_result_datain <= w_sys_tmp5711;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub21_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub21_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1c4: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub21_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h1b: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub28_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub28_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_u_addr <= $signed( w_sys_tmp2510[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_u_datain <= w_sys_tmp2513;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hcf: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub28_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub28_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp3131[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp3122[11:0] );

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp3125[11:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp3119[11:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp5249[11:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp5254[11:0] );

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub28_result_addr <= $signed( w_sys_tmp9828[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_sub28_result_datain <= w_sys_tmp3160;

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub28_result_datain <= r_sys_tmp2_float;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub28_result_datain <= w_sys_tmp5258;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub28_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub28_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub28_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub28_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub28_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h1c: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub29_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub29_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_u_addr <= $signed( w_sys_tmp2599[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_u_datain <= w_sys_tmp2602;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hd5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub29_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub29_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp3131[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp3122[11:0] );

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp3125[11:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp3119[11:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp5750[11:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp5755[11:0] );

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub29_result_addr <= $signed( w_sys_tmp9924[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub29_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub29_result_datain <= w_sys_tmp3171;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub29_result_datain <= w_sys_tmp5759;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub29_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub29_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub29_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1f9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub29_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub29_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h19: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub26_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub26_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_u_addr <= $signed( w_sys_tmp2332[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_u_datain <= w_sys_tmp2335;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc3: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub26_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub26_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp3131[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp3122[11:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp3125[11:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp3119[11:0] );

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp4252[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp4247[11:0] );

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub26_result_addr <= $signed( w_sys_tmp9636[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub26_result_datain <= w_sys_tmp3121;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub26_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub26_result_datain <= w_sys_tmp4256;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub26_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub26_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub26_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1e7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub26_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub26_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h8: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_u_addr <= $signed( w_sys_tmp839[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_u_datain <= w_sys_tmp842;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h53: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub09_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub09_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2963[11:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2951[11:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2957[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp2954[11:0] );

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3737[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3723[11:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3713[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp3708[11:0] );

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp8036[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub09_result_datain <= w_sys_tmp2959;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_datain <= w_sys_tmp3755;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub09_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub09_result_datain <= w_sys_tmp3717;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub09_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h177: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h1a: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub27_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub27_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_u_addr <= $signed( w_sys_tmp2421[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_u_datain <= w_sys_tmp2424;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hc9: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub27_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub27_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp3131[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp3122[11:0] );

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp3125[11:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp3119[11:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp4753[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp4748[11:0] );

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub27_result_addr <= $signed( w_sys_tmp9732[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub27_result_datain <= w_sys_tmp3149;

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub27_result_datain <= r_sys_tmp5_float;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub27_result_datain <= w_sys_tmp4757;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub27_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hf)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub27_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub27_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ed: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub27_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub27_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_u_addr <= $signed( w_sys_tmp762[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_u_datain <= w_sys_tmp765;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h4d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub08_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub08_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2960[11:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2951[11:0] );

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3236[11:0] );

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3212[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3222[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp3207[11:0] );

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp7959[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub08_result_datain <= w_sys_tmp2953;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub08_result_datain <= w_sys_tmp3254;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub08_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub08_result_datain <= w_sys_tmp3216;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub08_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h171: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h17: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub24_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub24_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_u_addr <= $signed( w_sys_tmp2166[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_u_datain <= w_sys_tmp2169;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hb7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub24_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub24_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp3128[11:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp3119[11:0] );

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp3250[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp3245[11:0] );

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp9463[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub24_result_datain <= w_sys_tmp3121;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub24_result_datain <= w_sys_tmp3254;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub24_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub24_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1db: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub24_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h18: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub25_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub25_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_u_addr <= $signed( w_sys_tmp2243[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_u_datain <= w_sys_tmp2246;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hbd: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub25_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub25_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp3131[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp3122[11:0] );

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp3125[11:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp3119[11:0] );

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp3746[11:0] );

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp3751[11:0] );

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub25_result_addr <= $signed( w_sys_tmp9540[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub25_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub25_result_datain <= w_sys_tmp3127;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub25_result_datain <= w_sys_tmp3755;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub25_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub25_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub25_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1e1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub25_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub25_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h15: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub22_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub22_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_u_addr <= $signed( w_sys_tmp1986[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_u_datain <= w_sys_tmp1989;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'ha6: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub22_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub22_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp3047[11:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp3035[11:0] );

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp3041[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp3038[11:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp6247[11:0] );

									end
									else
									if((r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h3b)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp6261[11:0] );

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp6237[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h34)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp6232[11:0] );

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp9268[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h19)) begin
										r_sub22_result_datain <= w_sys_tmp3098;

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub22_result_datain <= r_sys_tmp3_float;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub22_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub22_result_datain <= w_sys_tmp6212;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub22_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h14) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h1c) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h24) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h2c) || (r_sys_run_step==6'h33) || (r_sys_run_step==6'h34) || (r_sys_run_step==6'h3b)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub22_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ca: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub22_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h16: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub23_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub23_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_u_addr <= $signed( w_sys_tmp2075[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_u_datain <= w_sys_tmp2078;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hac: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub23_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub23_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp3041[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp3038[11:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp6738[11:0] );

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h3a)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp6748[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp6733[11:0] );

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp9364[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub23_result_datain <= w_sys_tmp3109;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h32)) begin
										r_sub23_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h39)) begin
										r_sub23_result_datain <= w_sys_tmp6713;

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub23_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'ha) || (r_sys_run_step==6'h2a)) begin
										r_sub23_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h22)) begin
										r_sub23_result_datain <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'h3a)) begin
										r_sub23_result_datain <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub23_result_datain <= r_sys_tmp2_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub23_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h11) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h21) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h29) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h31) || (r_sys_run_step==6'h32) || (r_sys_run_step==6'h39) || (r_sys_run_step==6'h3a)) begin
										r_sub23_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1d0: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub23_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h3: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_u_addr <= $signed( w_sys_tmp315[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_u_datain <= w_sys_tmp318;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h2a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub03_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub03_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2873[11:0] );

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2867[11:0] );

									end
									else
									if((r_sys_run_step==6'he)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2879[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2870[11:0] );

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4705[11:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp4720[11:0] );

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp7476[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'he)) begin
										r_sub03_result_datain <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==6'hd)) begin
										r_sub03_result_datain <= w_sys_tmp2897;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub03_result_datain <= w_sys_tmp4709;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hf)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'he)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub03_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h14e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h2: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_u_addr <= $signed( w_sys_tmp226[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_u_datain <= w_sys_tmp229;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h24: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub02_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub02_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2873[11:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2867[11:0] );

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2879[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2870[11:0] );

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp4219[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp4204[11:0] );

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp7380[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub02_result_datain <= w_sys_tmp2869;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub02_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub02_result_datain <= w_sys_tmp4208;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub02_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h148: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h1: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_u_addr <= $signed( w_sys_tmp137[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_u_datain <= w_sys_tmp140;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h1e: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub01_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub01_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2873[11:0] );

									end
									else
									if((r_sys_run_step==6'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2867[11:0] );

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2879[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2870[11:0] );

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3718[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp3703[11:0] );

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp7284[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h6)) begin
										r_sub01_result_datain <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==6'h5)) begin
										r_sub01_result_datain <= w_sys_tmp2875;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub01_result_datain <= w_sys_tmp3707;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub01_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h142: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_u_addr <= $signed( w_sys_tmp60[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_u_datain <= w_sys_tmp63;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h18: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub00_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub00_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2876[11:0] );

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2867[11:0] );

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3202[11:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp3217[11:0] );

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp7207[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_datain <= w_sys_tmp2869;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_datain <= w_sys_tmp3206;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub00_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h13c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h7: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_u_addr <= $signed( w_sys_tmp671[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_u_datain <= w_sys_tmp674;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h42: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub07_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub07_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2873[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2870[11:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp6724[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp6709[11:0] );

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp7860[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub07_result_datain <= w_sys_tmp2941;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub07_result_datain <= w_sys_tmp6713;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub07_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h166: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h6: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_u_addr <= $signed( w_sys_tmp582[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_u_datain <= w_sys_tmp585;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h3c: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub06_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub06_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h19)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2873[11:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2867[11:0] );

									end
									else
									if((r_sys_run_step==6'h1a)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2879[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2870[11:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp6208[11:0] );

									end
									else
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp6223[11:0] );

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp7764[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub06_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub06_result_datain <= w_sys_tmp2930;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub06_result_datain <= w_sys_tmp6212;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub06_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h160: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h5: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_u_addr <= $signed( w_sys_tmp493[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_u_datain <= w_sys_tmp496;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h36: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub05_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub05_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h15)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2873[11:0] );

									end
									else
									if((r_sys_run_step==6'h17)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2867[11:0] );

									end
									else
									if((r_sys_run_step==6'h16)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2879[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2870[11:0] );

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp5722[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp5707[11:0] );

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp7668[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h16)) begin
										r_sub05_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'h15)) begin
										r_sub05_result_datain <= w_sys_tmp2919;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub05_result_datain <= w_sys_tmp5711;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h17)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h15) || (r_sys_run_step==6'h16)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub05_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h15a: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h4: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_u_addr <= $signed( w_sys_tmp404[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_u_datain <= w_sys_tmp407;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h30: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub04_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub04_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h11)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2873[11:0] );

									end
									else
									if((r_sys_run_step==6'h13)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2867[11:0] );

									end
									else
									if((r_sys_run_step==6'h12)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2879[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2870[11:0] );

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp5221[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp5206[11:0] );

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp7572[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h12)) begin
										r_sub04_result_datain <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==6'h11)) begin
										r_sub04_result_datain <= w_sys_tmp2908;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_datain <= w_sys_tmp5210;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h13)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h11) || (r_sys_run_step==6'h12)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'h13) || (r_sys_run_step==6'h1b) || (r_sys_run_step==6'h23) || (r_sys_run_step==6'h2b) || (r_sys_run_step==6'h33)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'h12) || (r_sys_run_step==6'h1a) || (r_sys_run_step==6'h22) || (r_sys_run_step==6'h2a) || (r_sys_run_step==6'h32)) begin
										r_sub04_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h154: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h9: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_u_addr <= $signed( w_sys_tmp928[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_u_datain <= w_sys_tmp931;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h59: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub10_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub10_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'ha)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2963[11:0] );

									end
									else
									if((r_sys_run_step==6'hb)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2951[11:0] );

									end
									else
									if((r_sys_run_step==6'h9)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2957[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp2954[11:0] );

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4214[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4209[11:0] );

									end
									else
									if((r_sys_run_step==6'h6) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4224[11:0] );

									end
									else
									if((r_sys_run_step==6'h7) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h37)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp4238[11:0] );

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp8132[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sub10_result_datain <= w_sys_tmp2953;

									end
									else
									if((r_sys_run_step==6'ha)) begin
										r_sub10_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sub10_result_datain <= w_sys_tmp4218;

									end
									else
									if((r_sys_run_step==6'h6)) begin
										r_sub10_result_datain <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub10_result_datain <= w_sys_tmp4256;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'hb)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h9) || (r_sys_run_step==6'ha)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'hf) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h17) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h1f) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h27) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h2f) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h37)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h36)) begin
										r_sub10_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h17d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h1e: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub31_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub31_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_u_addr <= $signed( w_sys_tmp2777[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_u_datain <= w_sys_tmp2780;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he1: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub31_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub31_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp3122[11:0] );

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp3125[11:0] );

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp6752[11:0] );

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'he)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp6757[11:0] );

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub31_result_addr <= $signed( w_sys_tmp10116[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1d)) begin
										r_sub31_result_datain <= w_sys_tmp3193;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hc)) begin
										r_sub31_result_datain <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==6'h2)) begin
										r_sub31_result_datain <= w_sys_tmp6761;

									end
									else
									if((r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'ha)) begin
										r_sub31_result_datain <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==6'h8) || (r_sys_run_step==6'he)) begin
										r_sub31_result_datain <= r_sys_tmp1_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub31_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h1d)) begin
										r_sub31_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h3) || (r_sys_run_step==6'h5) || (r_sys_run_step==6'h7) || (r_sys_run_step==6'h9) || (r_sys_run_step==6'hb) || (r_sys_run_step==6'hd)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6) || (r_sys_run_step==6'h8) || (r_sys_run_step==6'ha) || (r_sys_run_step==6'hc) || (r_sys_run_step==6'he)) begin
										r_sub31_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h205: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub31_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub31_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h1d: begin
									if((r_sys_run_step==6'h1)) begin
										r_sub30_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub30_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_u_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_u_addr <= $signed( w_sys_tmp2688[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_u_datain <= w_sys_tmp2691;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_u_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hdb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h2<=r_sys_run_step && r_sys_run_step<=6'h8)) begin
										r_sub30_u_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_u_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub30_u_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_result_addr <= 12'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp3131[11:0] );

									end
									else
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp3122[11:0] );

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp3125[11:0] );

									end
									else
									if((r_sys_run_step==6'h1b)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp3119[11:0] );

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp6256[11:0] );

									end
									else
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp6251[11:0] );

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub30_result_addr <= $signed( w_sys_tmp10020[11:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h1a)) begin
										r_sub30_result_datain <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==6'h19)) begin
										r_sub30_result_datain <= w_sys_tmp3182;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub30_result_datain <= w_sys_tmp6260;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub30_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'he7: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h2: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h3: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h4: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h5: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h6: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h7: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h8: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h9: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'ha: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hb: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hc: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hd: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'he: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'hf: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h10: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h11: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h12: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h13: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h14: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h15: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h16: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h17: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h18: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h19: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1a: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1b: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1c: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1d: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

								6'h1e: begin
									if((r_sys_run_step==6'h0)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'h1b)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'h19) || (r_sys_run_step==6'h1a)) begin
										r_sub30_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h0) || (r_sys_run_step==6'he) || (r_sys_run_step==6'h16) || (r_sys_run_step==6'h1e) || (r_sys_run_step==6'h26) || (r_sys_run_step==6'h2e) || (r_sys_run_step==6'h36)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35) || (r_sys_run_step==6'h3d)) begin
										r_sub30_result_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						10'h1ff: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((6'h0<=r_sys_run_step && r_sys_run_step<=6'h6)) begin
										r_sub30_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						10'h207: begin
							r_sub30_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3)) begin
										r_sys_tmp0_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub26_result_dataout;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp0_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp0_float <= w_sub28_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5)) begin
										r_sys_tmp0_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp1_float <= w_sub27_result_dataout;

									end
								end

							endcase
						end

						10'h107: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp1_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp1_float <= w_sub29_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h5) || (r_sys_run_step==6'h8)) begin
										r_sys_tmp1_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub29_result_dataout;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp2_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						10'h119: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp2_float <= w_sub27_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sys_tmp2_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp3_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

						10'h10d: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp3_float <= w_sub25_result_dataout;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp3_float <= w_sub30_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'hb)) begin
										r_sys_tmp3_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub30_result_dataout;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						10'h11f: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub20_result_dataout;

									end
								end

							endcase
						end

						10'h125: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

						10'h12b: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp4_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'hd)) begin
										r_sys_tmp4_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'hef: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						10'hf5: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						10'hfb: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub20_result_dataout;

									end
								end

							endcase
						end

						10'h101: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2)) begin
										r_sys_tmp5_float <= w_sub28_result_dataout;

									end
								end

							endcase
						end

						10'h113: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'h10) || (r_sys_run_step==6'h18) || (r_sys_run_step==6'h20) || (r_sys_run_step==6'h28) || (r_sys_run_step==6'h30) || (r_sys_run_step==6'h38)) begin
										r_sys_tmp5_float <= w_sub26_result_dataout;

									end
								end

							endcase
						end

						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h9)) begin
										r_sys_tmp5_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h3) || (r_sys_run_step==6'h4) || (r_sys_run_step==6'h6)) begin
										r_sys_tmp6_float <= w_sub16_result_dataout;

									end
									else
									if((r_sys_run_step==6'hf)) begin
										r_sys_tmp6_float <= w_sub31_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						10'h131: begin

							case(r_sys_run_stage) 
								6'h0: begin
									if((r_sys_run_step==6'h7)) begin
										r_sys_tmp7_float <= w_sub16_result_dataout;

									end
									else
									if((r_sys_run_step==6'h2) || (r_sys_run_step==6'hd) || (r_sys_run_step==6'h15) || (r_sys_run_step==6'h1d) || (r_sys_run_step==6'h25) || (r_sys_run_step==6'h2d) || (r_sys_run_step==6'h35)) begin
										r_sys_tmp7_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
