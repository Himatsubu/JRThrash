/*
TimeStamp:	2016/6/1		8:13
*/


module P3(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg  signed [31:0] r_ip_DivInt_dividend_0;
	reg  signed [31:0] r_ip_DivInt_divisor_0;
	wire signed [31:0] w_ip_DivInt_quotient_0;
	wire signed [31:0] w_ip_DivInt_fractional_0;
	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 4:0] r_sys_run_stage;
	reg         [ 8:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 4:0] w_sys_run_stage_p1;
	wire        [ 8:0] w_sys_run_step_p1;
	wire signed [13:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [13:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [13:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [13:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [13:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [13:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [13:0] w_fld_V_3_addr_0;
	wire        [31:0] w_fld_V_3_datain_0;
	wire        [31:0] w_fld_V_3_dataout_0;
	wire               w_fld_V_3_r_w_0;
	wire               w_fld_V_3_ce_0;
	reg  signed [13:0] r_fld_V_3_addr_1;
	reg         [31:0] r_fld_V_3_datain_1;
	wire        [31:0] w_fld_V_3_dataout_1;
	reg                r_fld_V_3_r_w_1;
	wire               w_fld_V_3_ce_1;
	reg  signed [31:0] r_run_k_29;
	reg  signed [31:0] r_run_j_30;
	reg  signed [31:0] r_run_n_31;
	reg  signed [31:0] r_run_mx_32;
	reg  signed [31:0] r_run_my_33;
	reg         [31:0] r_run_dt_34;
	reg         [31:0] r_run_dx_35;
	reg         [31:0] r_run_dy_36;
	reg         [31:0] r_run_r1_37;
	reg         [31:0] r_run_r2_38;
	reg         [31:0] r_run_r3_39;
	reg         [31:0] r_run_r4_40;
	reg         [31:0] r_run_YY_41;
	reg  signed [31:0] r_run_kx_42;
	reg  signed [31:0] r_run_ky_43;
	reg  signed [31:0] r_run_nlast_44;
	reg  signed [31:0] r_run_copy0_j_45;
	reg  signed [31:0] r_run_copy1_j_46;
	reg  signed [31:0] r_run_copy2_j_47;
	reg  signed [31:0] r_run_copy0_j_48;
	reg                r_sub19_run_req;
	wire               w_sub19_run_busy;
	wire signed [13:0] w_sub19_T_addr;
	reg  signed [13:0] r_sub19_T_addr;
	wire        [31:0] w_sub19_T_datain;
	reg         [31:0] r_sub19_T_datain;
	wire        [31:0] w_sub19_T_dataout;
	wire               w_sub19_T_r_w;
	reg                r_sub19_T_r_w;
	wire signed [13:0] w_sub19_V_addr;
	reg  signed [13:0] r_sub19_V_addr;
	wire        [31:0] w_sub19_V_datain;
	reg         [31:0] r_sub19_V_datain;
	wire        [31:0] w_sub19_V_dataout;
	wire               w_sub19_V_r_w;
	reg                r_sub19_V_r_w;
	wire signed [13:0] w_sub19_U_addr;
	reg  signed [13:0] r_sub19_U_addr;
	wire        [31:0] w_sub19_U_datain;
	reg         [31:0] r_sub19_U_datain;
	wire        [31:0] w_sub19_U_dataout;
	wire               w_sub19_U_r_w;
	reg                r_sub19_U_r_w;
	wire signed [13:0] w_sub19_result_addr;
	reg  signed [13:0] r_sub19_result_addr;
	wire        [31:0] w_sub19_result_datain;
	reg         [31:0] r_sub19_result_datain;
	wire        [31:0] w_sub19_result_dataout;
	wire               w_sub19_result_r_w;
	reg                r_sub19_result_r_w;
	reg                r_sub09_run_req;
	wire               w_sub09_run_busy;
	wire signed [13:0] w_sub09_T_addr;
	reg  signed [13:0] r_sub09_T_addr;
	wire        [31:0] w_sub09_T_datain;
	reg         [31:0] r_sub09_T_datain;
	wire        [31:0] w_sub09_T_dataout;
	wire               w_sub09_T_r_w;
	reg                r_sub09_T_r_w;
	wire signed [13:0] w_sub09_V_addr;
	reg  signed [13:0] r_sub09_V_addr;
	wire        [31:0] w_sub09_V_datain;
	reg         [31:0] r_sub09_V_datain;
	wire        [31:0] w_sub09_V_dataout;
	wire               w_sub09_V_r_w;
	reg                r_sub09_V_r_w;
	wire signed [13:0] w_sub09_U_addr;
	reg  signed [13:0] r_sub09_U_addr;
	wire        [31:0] w_sub09_U_datain;
	reg         [31:0] r_sub09_U_datain;
	wire        [31:0] w_sub09_U_dataout;
	wire               w_sub09_U_r_w;
	reg                r_sub09_U_r_w;
	wire signed [13:0] w_sub09_result_addr;
	reg  signed [13:0] r_sub09_result_addr;
	wire        [31:0] w_sub09_result_datain;
	reg         [31:0] r_sub09_result_datain;
	wire        [31:0] w_sub09_result_dataout;
	wire               w_sub09_result_r_w;
	reg                r_sub09_result_r_w;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [13:0] w_sub08_T_addr;
	reg  signed [13:0] r_sub08_T_addr;
	wire        [31:0] w_sub08_T_datain;
	reg         [31:0] r_sub08_T_datain;
	wire        [31:0] w_sub08_T_dataout;
	wire               w_sub08_T_r_w;
	reg                r_sub08_T_r_w;
	wire signed [13:0] w_sub08_V_addr;
	reg  signed [13:0] r_sub08_V_addr;
	wire        [31:0] w_sub08_V_datain;
	reg         [31:0] r_sub08_V_datain;
	wire        [31:0] w_sub08_V_dataout;
	wire               w_sub08_V_r_w;
	reg                r_sub08_V_r_w;
	wire signed [13:0] w_sub08_U_addr;
	reg  signed [13:0] r_sub08_U_addr;
	wire        [31:0] w_sub08_U_datain;
	reg         [31:0] r_sub08_U_datain;
	wire        [31:0] w_sub08_U_dataout;
	wire               w_sub08_U_r_w;
	reg                r_sub08_U_r_w;
	wire signed [13:0] w_sub08_result_addr;
	reg  signed [13:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub24_run_req;
	wire               w_sub24_run_busy;
	wire signed [13:0] w_sub24_T_addr;
	reg  signed [13:0] r_sub24_T_addr;
	wire        [31:0] w_sub24_T_datain;
	reg         [31:0] r_sub24_T_datain;
	wire        [31:0] w_sub24_T_dataout;
	wire               w_sub24_T_r_w;
	reg                r_sub24_T_r_w;
	wire signed [13:0] w_sub24_V_addr;
	reg  signed [13:0] r_sub24_V_addr;
	wire        [31:0] w_sub24_V_datain;
	reg         [31:0] r_sub24_V_datain;
	wire        [31:0] w_sub24_V_dataout;
	wire               w_sub24_V_r_w;
	reg                r_sub24_V_r_w;
	wire signed [13:0] w_sub24_U_addr;
	reg  signed [13:0] r_sub24_U_addr;
	wire        [31:0] w_sub24_U_datain;
	reg         [31:0] r_sub24_U_datain;
	wire        [31:0] w_sub24_U_dataout;
	wire               w_sub24_U_r_w;
	reg                r_sub24_U_r_w;
	wire signed [13:0] w_sub24_result_addr;
	reg  signed [13:0] r_sub24_result_addr;
	wire        [31:0] w_sub24_result_datain;
	reg         [31:0] r_sub24_result_datain;
	wire        [31:0] w_sub24_result_dataout;
	wire               w_sub24_result_r_w;
	reg                r_sub24_result_r_w;
	reg                r_sub22_run_req;
	wire               w_sub22_run_busy;
	wire signed [13:0] w_sub22_T_addr;
	reg  signed [13:0] r_sub22_T_addr;
	wire        [31:0] w_sub22_T_datain;
	reg         [31:0] r_sub22_T_datain;
	wire        [31:0] w_sub22_T_dataout;
	wire               w_sub22_T_r_w;
	reg                r_sub22_T_r_w;
	wire signed [13:0] w_sub22_V_addr;
	reg  signed [13:0] r_sub22_V_addr;
	wire        [31:0] w_sub22_V_datain;
	reg         [31:0] r_sub22_V_datain;
	wire        [31:0] w_sub22_V_dataout;
	wire               w_sub22_V_r_w;
	reg                r_sub22_V_r_w;
	wire signed [13:0] w_sub22_U_addr;
	reg  signed [13:0] r_sub22_U_addr;
	wire        [31:0] w_sub22_U_datain;
	reg         [31:0] r_sub22_U_datain;
	wire        [31:0] w_sub22_U_dataout;
	wire               w_sub22_U_r_w;
	reg                r_sub22_U_r_w;
	wire signed [13:0] w_sub22_result_addr;
	reg  signed [13:0] r_sub22_result_addr;
	wire        [31:0] w_sub22_result_datain;
	reg         [31:0] r_sub22_result_datain;
	wire        [31:0] w_sub22_result_dataout;
	wire               w_sub22_result_r_w;
	reg                r_sub22_result_r_w;
	reg                r_sub23_run_req;
	wire               w_sub23_run_busy;
	wire signed [13:0] w_sub23_T_addr;
	reg  signed [13:0] r_sub23_T_addr;
	wire        [31:0] w_sub23_T_datain;
	reg         [31:0] r_sub23_T_datain;
	wire        [31:0] w_sub23_T_dataout;
	wire               w_sub23_T_r_w;
	reg                r_sub23_T_r_w;
	wire signed [13:0] w_sub23_V_addr;
	reg  signed [13:0] r_sub23_V_addr;
	wire        [31:0] w_sub23_V_datain;
	reg         [31:0] r_sub23_V_datain;
	wire        [31:0] w_sub23_V_dataout;
	wire               w_sub23_V_r_w;
	reg                r_sub23_V_r_w;
	wire signed [13:0] w_sub23_U_addr;
	reg  signed [13:0] r_sub23_U_addr;
	wire        [31:0] w_sub23_U_datain;
	reg         [31:0] r_sub23_U_datain;
	wire        [31:0] w_sub23_U_dataout;
	wire               w_sub23_U_r_w;
	reg                r_sub23_U_r_w;
	wire signed [13:0] w_sub23_result_addr;
	reg  signed [13:0] r_sub23_result_addr;
	wire        [31:0] w_sub23_result_datain;
	reg         [31:0] r_sub23_result_datain;
	wire        [31:0] w_sub23_result_dataout;
	wire               w_sub23_result_r_w;
	reg                r_sub23_result_r_w;
	reg                r_sub12_run_req;
	wire               w_sub12_run_busy;
	wire signed [13:0] w_sub12_T_addr;
	reg  signed [13:0] r_sub12_T_addr;
	wire        [31:0] w_sub12_T_datain;
	reg         [31:0] r_sub12_T_datain;
	wire        [31:0] w_sub12_T_dataout;
	wire               w_sub12_T_r_w;
	reg                r_sub12_T_r_w;
	wire signed [13:0] w_sub12_V_addr;
	reg  signed [13:0] r_sub12_V_addr;
	wire        [31:0] w_sub12_V_datain;
	reg         [31:0] r_sub12_V_datain;
	wire        [31:0] w_sub12_V_dataout;
	wire               w_sub12_V_r_w;
	reg                r_sub12_V_r_w;
	wire signed [13:0] w_sub12_U_addr;
	reg  signed [13:0] r_sub12_U_addr;
	wire        [31:0] w_sub12_U_datain;
	reg         [31:0] r_sub12_U_datain;
	wire        [31:0] w_sub12_U_dataout;
	wire               w_sub12_U_r_w;
	reg                r_sub12_U_r_w;
	wire signed [13:0] w_sub12_result_addr;
	reg  signed [13:0] r_sub12_result_addr;
	wire        [31:0] w_sub12_result_datain;
	reg         [31:0] r_sub12_result_datain;
	wire        [31:0] w_sub12_result_dataout;
	wire               w_sub12_result_r_w;
	reg                r_sub12_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [13:0] w_sub03_T_addr;
	reg  signed [13:0] r_sub03_T_addr;
	wire        [31:0] w_sub03_T_datain;
	reg         [31:0] r_sub03_T_datain;
	wire        [31:0] w_sub03_T_dataout;
	wire               w_sub03_T_r_w;
	reg                r_sub03_T_r_w;
	wire signed [13:0] w_sub03_V_addr;
	reg  signed [13:0] r_sub03_V_addr;
	wire        [31:0] w_sub03_V_datain;
	reg         [31:0] r_sub03_V_datain;
	wire        [31:0] w_sub03_V_dataout;
	wire               w_sub03_V_r_w;
	reg                r_sub03_V_r_w;
	wire signed [13:0] w_sub03_U_addr;
	reg  signed [13:0] r_sub03_U_addr;
	wire        [31:0] w_sub03_U_datain;
	reg         [31:0] r_sub03_U_datain;
	wire        [31:0] w_sub03_U_dataout;
	wire               w_sub03_U_r_w;
	reg                r_sub03_U_r_w;
	wire signed [13:0] w_sub03_result_addr;
	reg  signed [13:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [13:0] w_sub02_T_addr;
	reg  signed [13:0] r_sub02_T_addr;
	wire        [31:0] w_sub02_T_datain;
	reg         [31:0] r_sub02_T_datain;
	wire        [31:0] w_sub02_T_dataout;
	wire               w_sub02_T_r_w;
	reg                r_sub02_T_r_w;
	wire signed [13:0] w_sub02_V_addr;
	reg  signed [13:0] r_sub02_V_addr;
	wire        [31:0] w_sub02_V_datain;
	reg         [31:0] r_sub02_V_datain;
	wire        [31:0] w_sub02_V_dataout;
	wire               w_sub02_V_r_w;
	reg                r_sub02_V_r_w;
	wire signed [13:0] w_sub02_U_addr;
	reg  signed [13:0] r_sub02_U_addr;
	wire        [31:0] w_sub02_U_datain;
	reg         [31:0] r_sub02_U_datain;
	wire        [31:0] w_sub02_U_dataout;
	wire               w_sub02_U_r_w;
	reg                r_sub02_U_r_w;
	wire signed [13:0] w_sub02_result_addr;
	reg  signed [13:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub11_run_req;
	wire               w_sub11_run_busy;
	wire signed [13:0] w_sub11_T_addr;
	reg  signed [13:0] r_sub11_T_addr;
	wire        [31:0] w_sub11_T_datain;
	reg         [31:0] r_sub11_T_datain;
	wire        [31:0] w_sub11_T_dataout;
	wire               w_sub11_T_r_w;
	reg                r_sub11_T_r_w;
	wire signed [13:0] w_sub11_V_addr;
	reg  signed [13:0] r_sub11_V_addr;
	wire        [31:0] w_sub11_V_datain;
	reg         [31:0] r_sub11_V_datain;
	wire        [31:0] w_sub11_V_dataout;
	wire               w_sub11_V_r_w;
	reg                r_sub11_V_r_w;
	wire signed [13:0] w_sub11_U_addr;
	reg  signed [13:0] r_sub11_U_addr;
	wire        [31:0] w_sub11_U_datain;
	reg         [31:0] r_sub11_U_datain;
	wire        [31:0] w_sub11_U_dataout;
	wire               w_sub11_U_r_w;
	reg                r_sub11_U_r_w;
	wire signed [13:0] w_sub11_result_addr;
	reg  signed [13:0] r_sub11_result_addr;
	wire        [31:0] w_sub11_result_datain;
	reg         [31:0] r_sub11_result_datain;
	wire        [31:0] w_sub11_result_dataout;
	wire               w_sub11_result_r_w;
	reg                r_sub11_result_r_w;
	reg                r_sub14_run_req;
	wire               w_sub14_run_busy;
	wire signed [13:0] w_sub14_T_addr;
	reg  signed [13:0] r_sub14_T_addr;
	wire        [31:0] w_sub14_T_datain;
	reg         [31:0] r_sub14_T_datain;
	wire        [31:0] w_sub14_T_dataout;
	wire               w_sub14_T_r_w;
	reg                r_sub14_T_r_w;
	wire signed [13:0] w_sub14_V_addr;
	reg  signed [13:0] r_sub14_V_addr;
	wire        [31:0] w_sub14_V_datain;
	reg         [31:0] r_sub14_V_datain;
	wire        [31:0] w_sub14_V_dataout;
	wire               w_sub14_V_r_w;
	reg                r_sub14_V_r_w;
	wire signed [13:0] w_sub14_U_addr;
	reg  signed [13:0] r_sub14_U_addr;
	wire        [31:0] w_sub14_U_datain;
	reg         [31:0] r_sub14_U_datain;
	wire        [31:0] w_sub14_U_dataout;
	wire               w_sub14_U_r_w;
	reg                r_sub14_U_r_w;
	wire signed [13:0] w_sub14_result_addr;
	reg  signed [13:0] r_sub14_result_addr;
	wire        [31:0] w_sub14_result_datain;
	reg         [31:0] r_sub14_result_datain;
	wire        [31:0] w_sub14_result_dataout;
	wire               w_sub14_result_r_w;
	reg                r_sub14_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [13:0] w_sub01_T_addr;
	reg  signed [13:0] r_sub01_T_addr;
	wire        [31:0] w_sub01_T_datain;
	reg         [31:0] r_sub01_T_datain;
	wire        [31:0] w_sub01_T_dataout;
	wire               w_sub01_T_r_w;
	reg                r_sub01_T_r_w;
	wire signed [13:0] w_sub01_V_addr;
	reg  signed [13:0] r_sub01_V_addr;
	wire        [31:0] w_sub01_V_datain;
	reg         [31:0] r_sub01_V_datain;
	wire        [31:0] w_sub01_V_dataout;
	wire               w_sub01_V_r_w;
	reg                r_sub01_V_r_w;
	wire signed [13:0] w_sub01_U_addr;
	reg  signed [13:0] r_sub01_U_addr;
	wire        [31:0] w_sub01_U_datain;
	reg         [31:0] r_sub01_U_datain;
	wire        [31:0] w_sub01_U_dataout;
	wire               w_sub01_U_r_w;
	reg                r_sub01_U_r_w;
	wire signed [13:0] w_sub01_result_addr;
	reg  signed [13:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [13:0] w_sub00_T_addr;
	reg  signed [13:0] r_sub00_T_addr;
	wire        [31:0] w_sub00_T_datain;
	reg         [31:0] r_sub00_T_datain;
	wire        [31:0] w_sub00_T_dataout;
	wire               w_sub00_T_r_w;
	reg                r_sub00_T_r_w;
	wire signed [13:0] w_sub00_V_addr;
	reg  signed [13:0] r_sub00_V_addr;
	wire        [31:0] w_sub00_V_datain;
	reg         [31:0] r_sub00_V_datain;
	wire        [31:0] w_sub00_V_dataout;
	wire               w_sub00_V_r_w;
	reg                r_sub00_V_r_w;
	wire signed [13:0] w_sub00_U_addr;
	reg  signed [13:0] r_sub00_U_addr;
	wire        [31:0] w_sub00_U_datain;
	reg         [31:0] r_sub00_U_datain;
	wire        [31:0] w_sub00_U_dataout;
	wire               w_sub00_U_r_w;
	reg                r_sub00_U_r_w;
	wire signed [13:0] w_sub00_result_addr;
	reg  signed [13:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub13_run_req;
	wire               w_sub13_run_busy;
	wire signed [13:0] w_sub13_T_addr;
	reg  signed [13:0] r_sub13_T_addr;
	wire        [31:0] w_sub13_T_datain;
	reg         [31:0] r_sub13_T_datain;
	wire        [31:0] w_sub13_T_dataout;
	wire               w_sub13_T_r_w;
	reg                r_sub13_T_r_w;
	wire signed [13:0] w_sub13_V_addr;
	reg  signed [13:0] r_sub13_V_addr;
	wire        [31:0] w_sub13_V_datain;
	reg         [31:0] r_sub13_V_datain;
	wire        [31:0] w_sub13_V_dataout;
	wire               w_sub13_V_r_w;
	reg                r_sub13_V_r_w;
	wire signed [13:0] w_sub13_U_addr;
	reg  signed [13:0] r_sub13_U_addr;
	wire        [31:0] w_sub13_U_datain;
	reg         [31:0] r_sub13_U_datain;
	wire        [31:0] w_sub13_U_dataout;
	wire               w_sub13_U_r_w;
	reg                r_sub13_U_r_w;
	wire signed [13:0] w_sub13_result_addr;
	reg  signed [13:0] r_sub13_result_addr;
	wire        [31:0] w_sub13_result_datain;
	reg         [31:0] r_sub13_result_datain;
	wire        [31:0] w_sub13_result_dataout;
	wire               w_sub13_result_r_w;
	reg                r_sub13_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [13:0] w_sub07_T_addr;
	reg  signed [13:0] r_sub07_T_addr;
	wire        [31:0] w_sub07_T_datain;
	reg         [31:0] r_sub07_T_datain;
	wire        [31:0] w_sub07_T_dataout;
	wire               w_sub07_T_r_w;
	reg                r_sub07_T_r_w;
	wire signed [13:0] w_sub07_V_addr;
	reg  signed [13:0] r_sub07_V_addr;
	wire        [31:0] w_sub07_V_datain;
	reg         [31:0] r_sub07_V_datain;
	wire        [31:0] w_sub07_V_dataout;
	wire               w_sub07_V_r_w;
	reg                r_sub07_V_r_w;
	wire signed [13:0] w_sub07_U_addr;
	reg  signed [13:0] r_sub07_U_addr;
	wire        [31:0] w_sub07_U_datain;
	reg         [31:0] r_sub07_U_datain;
	wire        [31:0] w_sub07_U_dataout;
	wire               w_sub07_U_r_w;
	reg                r_sub07_U_r_w;
	wire signed [13:0] w_sub07_result_addr;
	reg  signed [13:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub16_run_req;
	wire               w_sub16_run_busy;
	wire signed [13:0] w_sub16_T_addr;
	reg  signed [13:0] r_sub16_T_addr;
	wire        [31:0] w_sub16_T_datain;
	reg         [31:0] r_sub16_T_datain;
	wire        [31:0] w_sub16_T_dataout;
	wire               w_sub16_T_r_w;
	reg                r_sub16_T_r_w;
	wire signed [13:0] w_sub16_V_addr;
	reg  signed [13:0] r_sub16_V_addr;
	wire        [31:0] w_sub16_V_datain;
	reg         [31:0] r_sub16_V_datain;
	wire        [31:0] w_sub16_V_dataout;
	wire               w_sub16_V_r_w;
	reg                r_sub16_V_r_w;
	wire signed [13:0] w_sub16_U_addr;
	reg  signed [13:0] r_sub16_U_addr;
	wire        [31:0] w_sub16_U_datain;
	reg         [31:0] r_sub16_U_datain;
	wire        [31:0] w_sub16_U_dataout;
	wire               w_sub16_U_r_w;
	reg                r_sub16_U_r_w;
	wire signed [13:0] w_sub16_result_addr;
	reg  signed [13:0] r_sub16_result_addr;
	wire        [31:0] w_sub16_result_datain;
	reg         [31:0] r_sub16_result_datain;
	wire        [31:0] w_sub16_result_dataout;
	wire               w_sub16_result_r_w;
	reg                r_sub16_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [13:0] w_sub06_T_addr;
	reg  signed [13:0] r_sub06_T_addr;
	wire        [31:0] w_sub06_T_datain;
	reg         [31:0] r_sub06_T_datain;
	wire        [31:0] w_sub06_T_dataout;
	wire               w_sub06_T_r_w;
	reg                r_sub06_T_r_w;
	wire signed [13:0] w_sub06_V_addr;
	reg  signed [13:0] r_sub06_V_addr;
	wire        [31:0] w_sub06_V_datain;
	reg         [31:0] r_sub06_V_datain;
	wire        [31:0] w_sub06_V_dataout;
	wire               w_sub06_V_r_w;
	reg                r_sub06_V_r_w;
	wire signed [13:0] w_sub06_U_addr;
	reg  signed [13:0] r_sub06_U_addr;
	wire        [31:0] w_sub06_U_datain;
	reg         [31:0] r_sub06_U_datain;
	wire        [31:0] w_sub06_U_dataout;
	wire               w_sub06_U_r_w;
	reg                r_sub06_U_r_w;
	wire signed [13:0] w_sub06_result_addr;
	reg  signed [13:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub15_run_req;
	wire               w_sub15_run_busy;
	wire signed [13:0] w_sub15_T_addr;
	reg  signed [13:0] r_sub15_T_addr;
	wire        [31:0] w_sub15_T_datain;
	reg         [31:0] r_sub15_T_datain;
	wire        [31:0] w_sub15_T_dataout;
	wire               w_sub15_T_r_w;
	reg                r_sub15_T_r_w;
	wire signed [13:0] w_sub15_V_addr;
	reg  signed [13:0] r_sub15_V_addr;
	wire        [31:0] w_sub15_V_datain;
	reg         [31:0] r_sub15_V_datain;
	wire        [31:0] w_sub15_V_dataout;
	wire               w_sub15_V_r_w;
	reg                r_sub15_V_r_w;
	wire signed [13:0] w_sub15_U_addr;
	reg  signed [13:0] r_sub15_U_addr;
	wire        [31:0] w_sub15_U_datain;
	reg         [31:0] r_sub15_U_datain;
	wire        [31:0] w_sub15_U_dataout;
	wire               w_sub15_U_r_w;
	reg                r_sub15_U_r_w;
	wire signed [13:0] w_sub15_result_addr;
	reg  signed [13:0] r_sub15_result_addr;
	wire        [31:0] w_sub15_result_datain;
	reg         [31:0] r_sub15_result_datain;
	wire        [31:0] w_sub15_result_dataout;
	wire               w_sub15_result_r_w;
	reg                r_sub15_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [13:0] w_sub05_T_addr;
	reg  signed [13:0] r_sub05_T_addr;
	wire        [31:0] w_sub05_T_datain;
	reg         [31:0] r_sub05_T_datain;
	wire        [31:0] w_sub05_T_dataout;
	wire               w_sub05_T_r_w;
	reg                r_sub05_T_r_w;
	wire signed [13:0] w_sub05_V_addr;
	reg  signed [13:0] r_sub05_V_addr;
	wire        [31:0] w_sub05_V_datain;
	reg         [31:0] r_sub05_V_datain;
	wire        [31:0] w_sub05_V_dataout;
	wire               w_sub05_V_r_w;
	reg                r_sub05_V_r_w;
	wire signed [13:0] w_sub05_U_addr;
	reg  signed [13:0] r_sub05_U_addr;
	wire        [31:0] w_sub05_U_datain;
	reg         [31:0] r_sub05_U_datain;
	wire        [31:0] w_sub05_U_dataout;
	wire               w_sub05_U_r_w;
	reg                r_sub05_U_r_w;
	wire signed [13:0] w_sub05_result_addr;
	reg  signed [13:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub18_run_req;
	wire               w_sub18_run_busy;
	wire signed [13:0] w_sub18_T_addr;
	reg  signed [13:0] r_sub18_T_addr;
	wire        [31:0] w_sub18_T_datain;
	reg         [31:0] r_sub18_T_datain;
	wire        [31:0] w_sub18_T_dataout;
	wire               w_sub18_T_r_w;
	reg                r_sub18_T_r_w;
	wire signed [13:0] w_sub18_V_addr;
	reg  signed [13:0] r_sub18_V_addr;
	wire        [31:0] w_sub18_V_datain;
	reg         [31:0] r_sub18_V_datain;
	wire        [31:0] w_sub18_V_dataout;
	wire               w_sub18_V_r_w;
	reg                r_sub18_V_r_w;
	wire signed [13:0] w_sub18_U_addr;
	reg  signed [13:0] r_sub18_U_addr;
	wire        [31:0] w_sub18_U_datain;
	reg         [31:0] r_sub18_U_datain;
	wire        [31:0] w_sub18_U_dataout;
	wire               w_sub18_U_r_w;
	reg                r_sub18_U_r_w;
	wire signed [13:0] w_sub18_result_addr;
	reg  signed [13:0] r_sub18_result_addr;
	wire        [31:0] w_sub18_result_datain;
	reg         [31:0] r_sub18_result_datain;
	wire        [31:0] w_sub18_result_dataout;
	wire               w_sub18_result_r_w;
	reg                r_sub18_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [13:0] w_sub04_T_addr;
	reg  signed [13:0] r_sub04_T_addr;
	wire        [31:0] w_sub04_T_datain;
	reg         [31:0] r_sub04_T_datain;
	wire        [31:0] w_sub04_T_dataout;
	wire               w_sub04_T_r_w;
	reg                r_sub04_T_r_w;
	wire signed [13:0] w_sub04_V_addr;
	reg  signed [13:0] r_sub04_V_addr;
	wire        [31:0] w_sub04_V_datain;
	reg         [31:0] r_sub04_V_datain;
	wire        [31:0] w_sub04_V_dataout;
	wire               w_sub04_V_r_w;
	reg                r_sub04_V_r_w;
	wire signed [13:0] w_sub04_U_addr;
	reg  signed [13:0] r_sub04_U_addr;
	wire        [31:0] w_sub04_U_datain;
	reg         [31:0] r_sub04_U_datain;
	wire        [31:0] w_sub04_U_dataout;
	wire               w_sub04_U_r_w;
	reg                r_sub04_U_r_w;
	wire signed [13:0] w_sub04_result_addr;
	reg  signed [13:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg                r_sub17_run_req;
	wire               w_sub17_run_busy;
	wire signed [13:0] w_sub17_T_addr;
	reg  signed [13:0] r_sub17_T_addr;
	wire        [31:0] w_sub17_T_datain;
	reg         [31:0] r_sub17_T_datain;
	wire        [31:0] w_sub17_T_dataout;
	wire               w_sub17_T_r_w;
	reg                r_sub17_T_r_w;
	wire signed [13:0] w_sub17_V_addr;
	reg  signed [13:0] r_sub17_V_addr;
	wire        [31:0] w_sub17_V_datain;
	reg         [31:0] r_sub17_V_datain;
	wire        [31:0] w_sub17_V_dataout;
	wire               w_sub17_V_r_w;
	reg                r_sub17_V_r_w;
	wire signed [13:0] w_sub17_U_addr;
	reg  signed [13:0] r_sub17_U_addr;
	wire        [31:0] w_sub17_U_datain;
	reg         [31:0] r_sub17_U_datain;
	wire        [31:0] w_sub17_U_dataout;
	wire               w_sub17_U_r_w;
	reg                r_sub17_U_r_w;
	wire signed [13:0] w_sub17_result_addr;
	reg  signed [13:0] r_sub17_result_addr;
	wire        [31:0] w_sub17_result_datain;
	reg         [31:0] r_sub17_result_datain;
	wire        [31:0] w_sub17_result_dataout;
	wire               w_sub17_result_r_w;
	reg                r_sub17_result_r_w;
	reg                r_sub10_run_req;
	wire               w_sub10_run_busy;
	wire signed [13:0] w_sub10_T_addr;
	reg  signed [13:0] r_sub10_T_addr;
	wire        [31:0] w_sub10_T_datain;
	reg         [31:0] r_sub10_T_datain;
	wire        [31:0] w_sub10_T_dataout;
	wire               w_sub10_T_r_w;
	reg                r_sub10_T_r_w;
	wire signed [13:0] w_sub10_V_addr;
	reg  signed [13:0] r_sub10_V_addr;
	wire        [31:0] w_sub10_V_datain;
	reg         [31:0] r_sub10_V_datain;
	wire        [31:0] w_sub10_V_dataout;
	wire               w_sub10_V_r_w;
	reg                r_sub10_V_r_w;
	wire signed [13:0] w_sub10_U_addr;
	reg  signed [13:0] r_sub10_U_addr;
	wire        [31:0] w_sub10_U_datain;
	reg         [31:0] r_sub10_U_datain;
	wire        [31:0] w_sub10_U_dataout;
	wire               w_sub10_U_r_w;
	reg                r_sub10_U_r_w;
	wire signed [13:0] w_sub10_result_addr;
	reg  signed [13:0] r_sub10_result_addr;
	wire        [31:0] w_sub10_result_datain;
	reg         [31:0] r_sub10_result_datain;
	wire        [31:0] w_sub10_result_dataout;
	wire               w_sub10_result_r_w;
	reg                r_sub10_result_r_w;
	reg                r_sub20_run_req;
	wire               w_sub20_run_busy;
	wire signed [13:0] w_sub20_T_addr;
	reg  signed [13:0] r_sub20_T_addr;
	wire        [31:0] w_sub20_T_datain;
	reg         [31:0] r_sub20_T_datain;
	wire        [31:0] w_sub20_T_dataout;
	wire               w_sub20_T_r_w;
	reg                r_sub20_T_r_w;
	wire signed [13:0] w_sub20_V_addr;
	reg  signed [13:0] r_sub20_V_addr;
	wire        [31:0] w_sub20_V_datain;
	reg         [31:0] r_sub20_V_datain;
	wire        [31:0] w_sub20_V_dataout;
	wire               w_sub20_V_r_w;
	reg                r_sub20_V_r_w;
	wire signed [13:0] w_sub20_U_addr;
	reg  signed [13:0] r_sub20_U_addr;
	wire        [31:0] w_sub20_U_datain;
	reg         [31:0] r_sub20_U_datain;
	wire        [31:0] w_sub20_U_dataout;
	wire               w_sub20_U_r_w;
	reg                r_sub20_U_r_w;
	wire signed [13:0] w_sub20_result_addr;
	reg  signed [13:0] r_sub20_result_addr;
	wire        [31:0] w_sub20_result_datain;
	reg         [31:0] r_sub20_result_datain;
	wire        [31:0] w_sub20_result_dataout;
	wire               w_sub20_result_r_w;
	reg                r_sub20_result_r_w;
	reg                r_sub21_run_req;
	wire               w_sub21_run_busy;
	wire signed [13:0] w_sub21_T_addr;
	reg  signed [13:0] r_sub21_T_addr;
	wire        [31:0] w_sub21_T_datain;
	reg         [31:0] r_sub21_T_datain;
	wire        [31:0] w_sub21_T_dataout;
	wire               w_sub21_T_r_w;
	reg                r_sub21_T_r_w;
	wire signed [13:0] w_sub21_V_addr;
	reg  signed [13:0] r_sub21_V_addr;
	wire        [31:0] w_sub21_V_datain;
	reg         [31:0] r_sub21_V_datain;
	wire        [31:0] w_sub21_V_dataout;
	wire               w_sub21_V_r_w;
	reg                r_sub21_V_r_w;
	wire signed [13:0] w_sub21_U_addr;
	reg  signed [13:0] r_sub21_U_addr;
	wire        [31:0] w_sub21_U_datain;
	reg         [31:0] r_sub21_U_datain;
	wire        [31:0] w_sub21_U_dataout;
	wire               w_sub21_U_r_w;
	reg                r_sub21_U_r_w;
	wire signed [13:0] w_sub21_result_addr;
	reg  signed [13:0] r_sub21_result_addr;
	wire        [31:0] w_sub21_result_datain;
	reg         [31:0] r_sub21_result_datain;
	wire        [31:0] w_sub21_result_dataout;
	wire               w_sub21_result_r_w;
	reg                r_sub21_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	reg         [31:0] r_sys_tmp48_float;
	reg         [31:0] r_sys_tmp49_float;
	reg         [31:0] r_sys_tmp50_float;
	reg         [31:0] r_sys_tmp51_float;
	reg         [31:0] r_sys_tmp52_float;
	reg         [31:0] r_sys_tmp53_float;
	reg         [31:0] r_sys_tmp54_float;
	reg         [31:0] r_sys_tmp55_float;
	reg         [31:0] r_sys_tmp56_float;
	reg         [31:0] r_sys_tmp57_float;
	reg         [31:0] r_sys_tmp58_float;
	reg         [31:0] r_sys_tmp59_float;
	reg         [31:0] r_sys_tmp60_float;
	reg         [31:0] r_sys_tmp61_float;
	reg         [31:0] r_sys_tmp62_float;
	reg         [31:0] r_sys_tmp63_float;
	reg         [31:0] r_sys_tmp64_float;
	reg         [31:0] r_sys_tmp65_float;
	reg         [31:0] r_sys_tmp66_float;
	reg         [31:0] r_sys_tmp67_float;
	reg         [31:0] r_sys_tmp68_float;
	reg         [31:0] r_sys_tmp69_float;
	reg         [31:0] r_sys_tmp70_float;
	reg         [31:0] r_sys_tmp71_float;
	reg         [31:0] r_sys_tmp72_float;
	reg         [31:0] r_sys_tmp73_float;
	reg         [31:0] r_sys_tmp74_float;
	reg         [31:0] r_sys_tmp75_float;
	reg         [31:0] r_sys_tmp76_float;
	reg         [31:0] r_sys_tmp77_float;
	reg         [31:0] r_sys_tmp78_float;
	reg         [31:0] r_sys_tmp79_float;
	reg         [31:0] r_sys_tmp80_float;
	reg         [31:0] r_sys_tmp81_float;
	reg         [31:0] r_sys_tmp82_float;
	reg         [31:0] r_sys_tmp83_float;
	reg         [31:0] r_sys_tmp84_float;
	reg         [31:0] r_sys_tmp85_float;
	reg         [31:0] r_sys_tmp86_float;
	reg         [31:0] r_sys_tmp87_float;
	reg         [31:0] r_sys_tmp88_float;
	reg         [31:0] r_sys_tmp89_float;
	reg         [31:0] r_sys_tmp90_float;
	reg         [31:0] r_sys_tmp91_float;
	reg         [31:0] r_sys_tmp92_float;
	reg         [31:0] r_sys_tmp93_float;
	reg         [31:0] r_sys_tmp94_float;
	reg         [31:0] r_sys_tmp95_float;
	reg         [31:0] r_sys_tmp96_float;
	reg         [31:0] r_sys_tmp97_float;
	reg         [31:0] r_sys_tmp98_float;
	reg         [31:0] r_sys_tmp99_float;
	reg         [31:0] r_sys_tmp100_float;
	reg         [31:0] r_sys_tmp101_float;
	reg         [31:0] r_sys_tmp102_float;
	reg         [31:0] r_sys_tmp103_float;
	reg         [31:0] r_sys_tmp104_float;
	reg         [31:0] r_sys_tmp105_float;
	reg         [31:0] r_sys_tmp106_float;
	reg         [31:0] r_sys_tmp107_float;
	reg         [31:0] r_sys_tmp108_float;
	reg         [31:0] r_sys_tmp109_float;
	reg         [31:0] r_sys_tmp110_float;
	reg         [31:0] r_sys_tmp111_float;
	reg         [31:0] r_sys_tmp112_float;
	reg         [31:0] r_sys_tmp113_float;
	reg         [31:0] r_sys_tmp114_float;
	reg         [31:0] r_sys_tmp115_float;
	reg         [31:0] r_sys_tmp116_float;
	reg         [31:0] r_sys_tmp117_float;
	reg         [31:0] r_sys_tmp118_float;
	reg         [31:0] r_sys_tmp119_float;
	reg         [31:0] r_sys_tmp120_float;
	reg         [31:0] r_sys_tmp121_float;
	reg         [31:0] r_sys_tmp122_float;
	reg         [31:0] r_sys_tmp123_float;
	reg         [31:0] r_sys_tmp124_float;
	reg         [31:0] r_sys_tmp125_float;
	reg         [31:0] r_sys_tmp126_float;
	reg         [31:0] r_sys_tmp127_float;
	reg         [31:0] r_sys_tmp128_float;
	reg         [31:0] r_sys_tmp129_float;
	reg         [31:0] r_sys_tmp130_float;
	reg         [31:0] r_sys_tmp131_float;
	reg         [31:0] r_sys_tmp132_float;
	reg         [31:0] r_sys_tmp133_float;
	reg         [31:0] r_sys_tmp134_float;
	reg         [31:0] r_sys_tmp135_float;
	reg         [31:0] r_sys_tmp136_float;
	reg         [31:0] r_sys_tmp137_float;
	reg         [31:0] r_sys_tmp138_float;
	reg         [31:0] r_sys_tmp139_float;
	reg         [31:0] r_sys_tmp140_float;
	reg         [31:0] r_sys_tmp141_float;
	reg         [31:0] r_sys_tmp142_float;
	reg         [31:0] r_sys_tmp143_float;
	reg         [31:0] r_sys_tmp144_float;
	reg         [31:0] r_sys_tmp145_float;
	reg         [31:0] r_sys_tmp146_float;
	reg         [31:0] r_sys_tmp147_float;
	reg         [31:0] r_sys_tmp148_float;
	reg         [31:0] r_sys_tmp149_float;
	reg         [31:0] r_sys_tmp150_float;
	reg         [31:0] r_sys_tmp151_float;
	reg         [31:0] r_sys_tmp152_float;
	reg         [31:0] r_sys_tmp153_float;
	reg         [31:0] r_sys_tmp154_float;
	reg         [31:0] r_sys_tmp155_float;
	reg         [31:0] r_sys_tmp156_float;
	reg         [31:0] r_sys_tmp157_float;
	reg         [31:0] r_sys_tmp158_float;
	reg         [31:0] r_sys_tmp159_float;
	reg         [31:0] r_sys_tmp160_float;
	reg         [31:0] r_sys_tmp161_float;
	reg         [31:0] r_sys_tmp162_float;
	reg         [31:0] r_sys_tmp163_float;
	reg         [31:0] r_sys_tmp164_float;
	reg         [31:0] r_sys_tmp165_float;
	reg         [31:0] r_sys_tmp166_float;
	reg         [31:0] r_sys_tmp167_float;
	reg         [31:0] r_sys_tmp168_float;
	reg         [31:0] r_sys_tmp169_float;
	reg         [31:0] r_sys_tmp170_float;
	reg         [31:0] r_sys_tmp171_float;
	reg         [31:0] r_sys_tmp172_float;
	reg         [31:0] r_sys_tmp173_float;
	reg         [31:0] r_sys_tmp174_float;
	reg         [31:0] r_sys_tmp175_float;
	reg         [31:0] r_sys_tmp176_float;
	reg         [31:0] r_sys_tmp177_float;
	reg         [31:0] r_sys_tmp178_float;
	reg         [31:0] r_sys_tmp179_float;
	reg         [31:0] r_sys_tmp180_float;
	reg         [31:0] r_sys_tmp181_float;
	reg         [31:0] r_sys_tmp182_float;
	reg         [31:0] r_sys_tmp183_float;
	reg         [31:0] r_sys_tmp184_float;
	reg         [31:0] r_sys_tmp185_float;
	reg         [31:0] r_sys_tmp186_float;
	reg         [31:0] r_sys_tmp187_float;
	reg         [31:0] r_sys_tmp188_float;
	reg         [31:0] r_sys_tmp189_float;
	reg         [31:0] r_sys_tmp190_float;
	reg         [31:0] r_sys_tmp191_float;
	reg         [31:0] r_sys_tmp192_float;
	reg         [31:0] r_sys_tmp193_float;
	reg         [31:0] r_sys_tmp194_float;
	reg         [31:0] r_sys_tmp195_float;
	reg         [31:0] r_sys_tmp196_float;
	reg         [31:0] r_sys_tmp197_float;
	reg         [31:0] r_sys_tmp198_float;
	reg         [31:0] r_sys_tmp199_float;
	reg         [31:0] r_sys_tmp200_float;
	reg         [31:0] r_sys_tmp201_float;
	reg         [31:0] r_sys_tmp202_float;
	reg         [31:0] r_sys_tmp203_float;
	reg         [31:0] r_sys_tmp204_float;
	reg         [31:0] r_sys_tmp205_float;
	reg         [31:0] r_sys_tmp206_float;
	reg         [31:0] r_sys_tmp207_float;
	reg         [31:0] r_sys_tmp208_float;
	reg         [31:0] r_sys_tmp209_float;
	reg         [31:0] r_sys_tmp210_float;
	reg         [31:0] r_sys_tmp211_float;
	reg         [31:0] r_sys_tmp212_float;
	reg         [31:0] r_sys_tmp213_float;
	reg         [31:0] r_sys_tmp214_float;
	reg         [31:0] r_sys_tmp215_float;
	reg         [31:0] r_sys_tmp216_float;
	reg         [31:0] r_sys_tmp217_float;
	reg         [31:0] r_sys_tmp218_float;
	reg         [31:0] r_sys_tmp219_float;
	reg         [31:0] r_sys_tmp220_float;
	reg         [31:0] r_sys_tmp221_float;
	reg         [31:0] r_sys_tmp222_float;
	reg         [31:0] r_sys_tmp223_float;
	reg         [31:0] r_sys_tmp224_float;
	reg         [31:0] r_sys_tmp225_float;
	reg         [31:0] r_sys_tmp226_float;
	reg         [31:0] r_sys_tmp227_float;
	reg         [31:0] r_sys_tmp228_float;
	reg         [31:0] r_sys_tmp229_float;
	reg         [31:0] r_sys_tmp230_float;
	reg         [31:0] r_sys_tmp231_float;
	reg         [31:0] r_sys_tmp232_float;
	reg         [31:0] r_sys_tmp233_float;
	reg         [31:0] r_sys_tmp234_float;
	reg         [31:0] r_sys_tmp235_float;
	reg         [31:0] r_sys_tmp236_float;
	reg         [31:0] r_sys_tmp237_float;
	reg         [31:0] r_sys_tmp238_float;
	reg         [31:0] r_sys_tmp239_float;
	reg         [31:0] r_sys_tmp240_float;
	reg         [31:0] r_sys_tmp241_float;
	reg         [31:0] r_sys_tmp242_float;
	reg         [31:0] r_sys_tmp243_float;
	reg         [31:0] r_sys_tmp244_float;
	reg         [31:0] r_sys_tmp245_float;
	reg         [31:0] r_sys_tmp246_float;
	reg         [31:0] r_sys_tmp247_float;
	reg         [31:0] r_sys_tmp248_float;
	reg         [31:0] r_sys_tmp249_float;
	reg         [31:0] r_sys_tmp250_float;
	reg         [31:0] r_sys_tmp251_float;
	reg         [31:0] r_sys_tmp252_float;
	reg         [31:0] r_sys_tmp253_float;
	reg         [31:0] r_sys_tmp254_float;
	reg         [31:0] r_sys_tmp255_float;
	reg         [31:0] r_sys_tmp256_float;
	reg         [31:0] r_sys_tmp257_float;
	reg         [31:0] r_sys_tmp258_float;
	reg         [31:0] r_sys_tmp259_float;
	reg         [31:0] r_sys_tmp260_float;
	reg         [31:0] r_sys_tmp261_float;
	reg         [31:0] r_sys_tmp262_float;
	reg         [31:0] r_sys_tmp263_float;
	reg         [31:0] r_sys_tmp264_float;
	reg         [31:0] r_sys_tmp265_float;
	reg         [31:0] r_sys_tmp266_float;
	reg         [31:0] r_sys_tmp267_float;
	reg         [31:0] r_sys_tmp268_float;
	reg         [31:0] r_sys_tmp269_float;
	reg         [31:0] r_sys_tmp270_float;
	reg         [31:0] r_sys_tmp271_float;
	reg         [31:0] r_sys_tmp272_float;
	reg         [31:0] r_sys_tmp273_float;
	reg         [31:0] r_sys_tmp274_float;
	reg         [31:0] r_sys_tmp275_float;
	reg         [31:0] r_sys_tmp276_float;
	reg         [31:0] r_sys_tmp277_float;
	reg         [31:0] r_sys_tmp278_float;
	reg         [31:0] r_sys_tmp279_float;
	reg         [31:0] r_sys_tmp280_float;
	reg         [31:0] r_sys_tmp281_float;
	reg         [31:0] r_sys_tmp282_float;
	reg         [31:0] r_sys_tmp283_float;
	reg         [31:0] r_sys_tmp284_float;
	reg         [31:0] r_sys_tmp285_float;
	reg         [31:0] r_sys_tmp286_float;
	reg         [31:0] r_sys_tmp287_float;
	reg         [31:0] r_sys_tmp288_float;
	reg         [31:0] r_sys_tmp289_float;
	reg         [31:0] r_sys_tmp290_float;
	reg         [31:0] r_sys_tmp291_float;
	reg         [31:0] r_sys_tmp292_float;
	reg         [31:0] r_sys_tmp293_float;
	reg         [31:0] r_sys_tmp294_float;
	reg         [31:0] r_sys_tmp295_float;
	reg         [31:0] r_sys_tmp296_float;
	reg         [31:0] r_sys_tmp297_float;
	reg         [31:0] r_sys_tmp298_float;
	reg         [31:0] r_sys_tmp299_float;
	reg         [31:0] r_sys_tmp300_float;
	reg         [31:0] r_sys_tmp301_float;
	reg         [31:0] r_sys_tmp302_float;
	reg         [31:0] r_sys_tmp303_float;
	reg         [31:0] r_sys_tmp304_float;
	reg         [31:0] r_sys_tmp305_float;
	reg         [31:0] r_sys_tmp306_float;
	reg         [31:0] r_sys_tmp307_float;
	reg         [31:0] r_sys_tmp308_float;
	reg         [31:0] r_sys_tmp309_float;
	reg         [31:0] r_sys_tmp310_float;
	reg         [31:0] r_sys_tmp311_float;
	reg         [31:0] r_sys_tmp312_float;
	reg         [31:0] r_sys_tmp313_float;
	reg         [31:0] r_sys_tmp314_float;
	reg         [31:0] r_sys_tmp315_float;
	reg         [31:0] r_sys_tmp316_float;
	reg         [31:0] r_sys_tmp317_float;
	reg         [31:0] r_sys_tmp318_float;
	reg         [31:0] r_sys_tmp319_float;
	reg         [31:0] r_sys_tmp320_float;
	reg         [31:0] r_sys_tmp321_float;
	reg         [31:0] r_sys_tmp322_float;
	reg         [31:0] r_sys_tmp323_float;
	reg         [31:0] r_sys_tmp324_float;
	reg         [31:0] r_sys_tmp325_float;
	reg         [31:0] r_sys_tmp326_float;
	reg         [31:0] r_sys_tmp327_float;
	reg         [31:0] r_sys_tmp328_float;
	reg         [31:0] r_sys_tmp329_float;
	reg         [31:0] r_sys_tmp330_float;
	reg         [31:0] r_sys_tmp331_float;
	reg         [31:0] r_sys_tmp332_float;
	reg         [31:0] r_sys_tmp333_float;
	reg         [31:0] r_sys_tmp334_float;
	reg         [31:0] r_sys_tmp335_float;
	reg         [31:0] r_sys_tmp336_float;
	reg         [31:0] r_sys_tmp337_float;
	reg         [31:0] r_sys_tmp338_float;
	reg         [31:0] r_sys_tmp339_float;
	reg         [31:0] r_sys_tmp340_float;
	reg         [31:0] r_sys_tmp341_float;
	reg         [31:0] r_sys_tmp342_float;
	reg         [31:0] r_sys_tmp343_float;
	reg         [31:0] r_sys_tmp344_float;
	reg         [31:0] r_sys_tmp345_float;
	reg         [31:0] r_sys_tmp346_float;
	reg         [31:0] r_sys_tmp347_float;
	reg         [31:0] r_sys_tmp348_float;
	reg         [31:0] r_sys_tmp349_float;
	reg         [31:0] r_sys_tmp350_float;
	reg         [31:0] r_sys_tmp351_float;
	reg         [31:0] r_sys_tmp352_float;
	reg         [31:0] r_sys_tmp353_float;
	reg         [31:0] r_sys_tmp354_float;
	reg         [31:0] r_sys_tmp355_float;
	reg         [31:0] r_sys_tmp356_float;
	reg         [31:0] r_sys_tmp357_float;
	reg         [31:0] r_sys_tmp358_float;
	reg         [31:0] r_sys_tmp359_float;
	reg         [31:0] r_sys_tmp360_float;
	reg         [31:0] r_sys_tmp361_float;
	reg         [31:0] r_sys_tmp362_float;
	reg         [31:0] r_sys_tmp363_float;
	reg         [31:0] r_sys_tmp364_float;
	reg         [31:0] r_sys_tmp365_float;
	reg         [31:0] r_sys_tmp366_float;
	reg         [31:0] r_sys_tmp367_float;
	reg         [31:0] r_sys_tmp368_float;
	reg         [31:0] r_sys_tmp369_float;
	reg         [31:0] r_sys_tmp370_float;
	reg         [31:0] r_sys_tmp371_float;
	reg         [31:0] r_sys_tmp372_float;
	reg         [31:0] r_sys_tmp373_float;
	reg         [31:0] r_sys_tmp374_float;
	reg         [31:0] r_sys_tmp375_float;
	reg         [31:0] r_sys_tmp376_float;
	reg         [31:0] r_sys_tmp377_float;
	reg         [31:0] r_sys_tmp378_float;
	reg         [31:0] r_sys_tmp379_float;
	reg         [31:0] r_sys_tmp380_float;
	reg         [31:0] r_sys_tmp381_float;
	reg         [31:0] r_sys_tmp382_float;
	reg         [31:0] r_sys_tmp383_float;
	reg         [31:0] r_sys_tmp384_float;
	reg         [31:0] r_sys_tmp385_float;
	reg         [31:0] r_sys_tmp386_float;
	reg         [31:0] r_sys_tmp387_float;
	reg         [31:0] r_sys_tmp388_float;
	reg         [31:0] r_sys_tmp389_float;
	reg         [31:0] r_sys_tmp390_float;
	reg         [31:0] r_sys_tmp391_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire        [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire               w_sys_tmp12;
	wire               w_sys_tmp13;
	wire signed [31:0] w_sys_tmp14;
	wire               w_sys_tmp15;
	wire               w_sys_tmp16;
	wire        [31:0] w_sys_tmp18;
	wire        [31:0] w_sys_tmp19;
	wire signed [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp22;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire        [31:0] w_sys_tmp25;
	wire signed [31:0] w_sys_tmp27;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp32;
	wire signed [31:0] w_sys_tmp33;
	wire        [31:0] w_sys_tmp36;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire signed [31:0] w_sys_tmp41;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp45;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire        [31:0] w_sys_tmp128;
	wire        [31:0] w_sys_tmp157;
	wire        [31:0] w_sys_tmp185;
	wire        [31:0] w_sys_tmp213;
	wire        [31:0] w_sys_tmp269;
	wire        [31:0] w_sys_tmp297;
	wire               w_sys_tmp588;
	wire               w_sys_tmp589;
	wire signed [31:0] w_sys_tmp590;
	wire signed [31:0] w_sys_tmp593;
	wire signed [31:0] w_sys_tmp594;
	wire        [31:0] w_sys_tmp595;
	wire        [31:0] w_sys_tmp601;
	wire signed [31:0] w_sys_tmp605;
	wire signed [31:0] w_sys_tmp606;
	wire signed [31:0] w_sys_tmp617;
	wire signed [31:0] w_sys_tmp618;
	wire signed [31:0] w_sys_tmp629;
	wire signed [31:0] w_sys_tmp630;
	wire signed [31:0] w_sys_tmp641;
	wire signed [31:0] w_sys_tmp642;
	wire signed [31:0] w_sys_tmp653;
	wire signed [31:0] w_sys_tmp654;
	wire signed [31:0] w_sys_tmp665;
	wire signed [31:0] w_sys_tmp666;
	wire signed [31:0] w_sys_tmp677;
	wire signed [31:0] w_sys_tmp678;
	wire signed [31:0] w_sys_tmp689;
	wire signed [31:0] w_sys_tmp690;
	wire signed [31:0] w_sys_tmp701;
	wire signed [31:0] w_sys_tmp702;
	wire signed [31:0] w_sys_tmp713;
	wire signed [31:0] w_sys_tmp714;
	wire signed [31:0] w_sys_tmp725;
	wire signed [31:0] w_sys_tmp726;
	wire signed [31:0] w_sys_tmp737;
	wire signed [31:0] w_sys_tmp738;
	wire signed [31:0] w_sys_tmp749;
	wire signed [31:0] w_sys_tmp750;
	wire signed [31:0] w_sys_tmp761;
	wire signed [31:0] w_sys_tmp762;
	wire signed [31:0] w_sys_tmp773;
	wire signed [31:0] w_sys_tmp774;
	wire signed [31:0] w_sys_tmp785;
	wire signed [31:0] w_sys_tmp786;
	wire signed [31:0] w_sys_tmp797;
	wire signed [31:0] w_sys_tmp798;
	wire signed [31:0] w_sys_tmp809;
	wire signed [31:0] w_sys_tmp810;
	wire signed [31:0] w_sys_tmp821;
	wire signed [31:0] w_sys_tmp822;
	wire signed [31:0] w_sys_tmp833;
	wire signed [31:0] w_sys_tmp834;
	wire signed [31:0] w_sys_tmp845;
	wire signed [31:0] w_sys_tmp846;
	wire signed [31:0] w_sys_tmp881;
	wire signed [31:0] w_sys_tmp882;
	wire signed [31:0] w_sys_tmp893;
	wire signed [31:0] w_sys_tmp894;
	wire signed [31:0] w_sys_tmp905;
	wire signed [31:0] w_sys_tmp906;
	wire signed [31:0] w_sys_tmp917;
	wire signed [31:0] w_sys_tmp918;
	wire signed [31:0] w_sys_tmp929;
	wire signed [31:0] w_sys_tmp930;
	wire signed [31:0] w_sys_tmp941;
	wire signed [31:0] w_sys_tmp942;
	wire signed [31:0] w_sys_tmp953;
	wire signed [31:0] w_sys_tmp954;
	wire signed [31:0] w_sys_tmp965;
	wire signed [31:0] w_sys_tmp966;
	wire signed [31:0] w_sys_tmp977;
	wire signed [31:0] w_sys_tmp978;
	wire signed [31:0] w_sys_tmp989;
	wire signed [31:0] w_sys_tmp990;
	wire signed [31:0] w_sys_tmp1001;
	wire signed [31:0] w_sys_tmp1002;
	wire signed [31:0] w_sys_tmp1013;
	wire signed [31:0] w_sys_tmp1014;
	wire signed [31:0] w_sys_tmp1025;
	wire signed [31:0] w_sys_tmp1026;
	wire signed [31:0] w_sys_tmp1037;
	wire signed [31:0] w_sys_tmp1038;
	wire signed [31:0] w_sys_tmp1049;
	wire signed [31:0] w_sys_tmp1050;
	wire signed [31:0] w_sys_tmp1061;
	wire signed [31:0] w_sys_tmp1062;
	wire signed [31:0] w_sys_tmp1073;
	wire signed [31:0] w_sys_tmp1074;
	wire signed [31:0] w_sys_tmp1085;
	wire signed [31:0] w_sys_tmp1086;
	wire signed [31:0] w_sys_tmp1097;
	wire signed [31:0] w_sys_tmp1098;
	wire signed [31:0] w_sys_tmp1109;
	wire signed [31:0] w_sys_tmp1110;
	wire signed [31:0] w_sys_tmp1145;
	wire signed [31:0] w_sys_tmp1146;
	wire signed [31:0] w_sys_tmp1157;
	wire signed [31:0] w_sys_tmp1158;
	wire signed [31:0] w_sys_tmp1169;
	wire signed [31:0] w_sys_tmp1170;
	wire signed [31:0] w_sys_tmp1181;
	wire signed [31:0] w_sys_tmp1182;
	wire signed [31:0] w_sys_tmp1193;
	wire signed [31:0] w_sys_tmp1194;
	wire signed [31:0] w_sys_tmp1205;
	wire signed [31:0] w_sys_tmp1206;
	wire signed [31:0] w_sys_tmp1217;
	wire signed [31:0] w_sys_tmp1218;
	wire signed [31:0] w_sys_tmp1229;
	wire signed [31:0] w_sys_tmp1230;
	wire signed [31:0] w_sys_tmp1241;
	wire signed [31:0] w_sys_tmp1242;
	wire signed [31:0] w_sys_tmp1253;
	wire signed [31:0] w_sys_tmp1254;
	wire signed [31:0] w_sys_tmp1265;
	wire signed [31:0] w_sys_tmp1266;
	wire signed [31:0] w_sys_tmp1277;
	wire signed [31:0] w_sys_tmp1278;
	wire signed [31:0] w_sys_tmp1289;
	wire signed [31:0] w_sys_tmp1290;
	wire signed [31:0] w_sys_tmp1301;
	wire signed [31:0] w_sys_tmp1302;
	wire signed [31:0] w_sys_tmp1313;
	wire signed [31:0] w_sys_tmp1314;
	wire signed [31:0] w_sys_tmp1325;
	wire signed [31:0] w_sys_tmp1326;
	wire signed [31:0] w_sys_tmp1337;
	wire signed [31:0] w_sys_tmp1338;
	wire signed [31:0] w_sys_tmp1349;
	wire signed [31:0] w_sys_tmp1350;
	wire signed [31:0] w_sys_tmp1361;
	wire signed [31:0] w_sys_tmp1362;
	wire signed [31:0] w_sys_tmp1385;
	wire signed [31:0] w_sys_tmp1386;
	wire signed [31:0] w_sys_tmp1397;
	wire signed [31:0] w_sys_tmp1398;
	wire signed [31:0] w_sys_tmp1409;
	wire signed [31:0] w_sys_tmp1410;
	wire signed [31:0] w_sys_tmp1421;
	wire signed [31:0] w_sys_tmp1422;
	wire signed [31:0] w_sys_tmp1433;
	wire signed [31:0] w_sys_tmp1434;
	wire signed [31:0] w_sys_tmp1445;
	wire signed [31:0] w_sys_tmp1446;
	wire signed [31:0] w_sys_tmp1457;
	wire signed [31:0] w_sys_tmp1458;
	wire signed [31:0] w_sys_tmp1469;
	wire signed [31:0] w_sys_tmp1470;
	wire signed [31:0] w_sys_tmp1481;
	wire signed [31:0] w_sys_tmp1482;
	wire signed [31:0] w_sys_tmp1493;
	wire signed [31:0] w_sys_tmp1494;
	wire signed [31:0] w_sys_tmp1505;
	wire signed [31:0] w_sys_tmp1506;
	wire signed [31:0] w_sys_tmp1517;
	wire signed [31:0] w_sys_tmp1518;
	wire signed [31:0] w_sys_tmp1529;
	wire signed [31:0] w_sys_tmp1530;
	wire signed [31:0] w_sys_tmp1541;
	wire signed [31:0] w_sys_tmp1542;
	wire signed [31:0] w_sys_tmp1553;
	wire signed [31:0] w_sys_tmp1554;
	wire signed [31:0] w_sys_tmp1565;
	wire signed [31:0] w_sys_tmp1566;
	wire signed [31:0] w_sys_tmp1577;
	wire signed [31:0] w_sys_tmp1578;
	wire signed [31:0] w_sys_tmp1589;
	wire signed [31:0] w_sys_tmp1590;
	wire signed [31:0] w_sys_tmp1601;
	wire signed [31:0] w_sys_tmp1602;
	wire signed [31:0] w_sys_tmp1613;
	wire signed [31:0] w_sys_tmp1614;
	wire signed [31:0] w_sys_tmp1625;
	wire signed [31:0] w_sys_tmp1626;
	wire signed [31:0] w_sys_tmp1661;
	wire signed [31:0] w_sys_tmp1662;
	wire signed [31:0] w_sys_tmp1673;
	wire signed [31:0] w_sys_tmp1674;
	wire signed [31:0] w_sys_tmp1685;
	wire signed [31:0] w_sys_tmp1686;
	wire signed [31:0] w_sys_tmp1697;
	wire signed [31:0] w_sys_tmp1698;
	wire signed [31:0] w_sys_tmp1709;
	wire signed [31:0] w_sys_tmp1710;
	wire signed [31:0] w_sys_tmp1721;
	wire signed [31:0] w_sys_tmp1722;
	wire signed [31:0] w_sys_tmp1733;
	wire signed [31:0] w_sys_tmp1734;
	wire signed [31:0] w_sys_tmp1745;
	wire signed [31:0] w_sys_tmp1746;
	wire signed [31:0] w_sys_tmp1757;
	wire signed [31:0] w_sys_tmp1758;
	wire signed [31:0] w_sys_tmp1769;
	wire signed [31:0] w_sys_tmp1770;
	wire signed [31:0] w_sys_tmp1781;
	wire signed [31:0] w_sys_tmp1782;
	wire signed [31:0] w_sys_tmp1793;
	wire signed [31:0] w_sys_tmp1794;
	wire signed [31:0] w_sys_tmp1805;
	wire signed [31:0] w_sys_tmp1806;
	wire signed [31:0] w_sys_tmp1817;
	wire signed [31:0] w_sys_tmp1818;
	wire signed [31:0] w_sys_tmp1829;
	wire signed [31:0] w_sys_tmp1830;
	wire signed [31:0] w_sys_tmp1841;
	wire signed [31:0] w_sys_tmp1842;
	wire signed [31:0] w_sys_tmp1853;
	wire signed [31:0] w_sys_tmp1854;
	wire signed [31:0] w_sys_tmp1865;
	wire signed [31:0] w_sys_tmp1866;
	wire signed [31:0] w_sys_tmp1877;
	wire signed [31:0] w_sys_tmp1878;
	wire signed [31:0] w_sys_tmp1889;
	wire signed [31:0] w_sys_tmp1890;
	wire signed [31:0] w_sys_tmp1901;
	wire signed [31:0] w_sys_tmp1902;
	wire signed [31:0] w_sys_tmp1913;
	wire signed [31:0] w_sys_tmp1914;
	wire signed [31:0] w_sys_tmp1925;
	wire signed [31:0] w_sys_tmp1926;
	wire signed [31:0] w_sys_tmp1937;
	wire signed [31:0] w_sys_tmp1938;
	wire signed [31:0] w_sys_tmp1949;
	wire signed [31:0] w_sys_tmp1950;
	wire signed [31:0] w_sys_tmp1961;
	wire signed [31:0] w_sys_tmp1962;
	wire signed [31:0] w_sys_tmp1973;
	wire signed [31:0] w_sys_tmp1974;
	wire signed [31:0] w_sys_tmp1985;
	wire signed [31:0] w_sys_tmp1986;
	wire signed [31:0] w_sys_tmp1997;
	wire signed [31:0] w_sys_tmp1998;
	wire signed [31:0] w_sys_tmp2009;
	wire signed [31:0] w_sys_tmp2010;
	wire signed [31:0] w_sys_tmp2021;
	wire signed [31:0] w_sys_tmp2022;
	wire signed [31:0] w_sys_tmp2033;
	wire signed [31:0] w_sys_tmp2034;
	wire signed [31:0] w_sys_tmp2045;
	wire signed [31:0] w_sys_tmp2046;
	wire signed [31:0] w_sys_tmp2057;
	wire signed [31:0] w_sys_tmp2058;
	wire signed [31:0] w_sys_tmp2069;
	wire signed [31:0] w_sys_tmp2070;
	wire signed [31:0] w_sys_tmp2081;
	wire signed [31:0] w_sys_tmp2082;
	wire signed [31:0] w_sys_tmp2093;
	wire signed [31:0] w_sys_tmp2094;
	wire signed [31:0] w_sys_tmp2105;
	wire signed [31:0] w_sys_tmp2106;
	wire signed [31:0] w_sys_tmp2117;
	wire signed [31:0] w_sys_tmp2118;
	wire signed [31:0] w_sys_tmp2129;
	wire signed [31:0] w_sys_tmp2130;
	wire signed [31:0] w_sys_tmp2153;
	wire signed [31:0] w_sys_tmp2154;
	wire signed [31:0] w_sys_tmp2165;
	wire signed [31:0] w_sys_tmp2166;
	wire signed [31:0] w_sys_tmp2177;
	wire signed [31:0] w_sys_tmp2178;
	wire signed [31:0] w_sys_tmp2189;
	wire signed [31:0] w_sys_tmp2190;
	wire signed [31:0] w_sys_tmp2201;
	wire signed [31:0] w_sys_tmp2202;
	wire signed [31:0] w_sys_tmp2213;
	wire signed [31:0] w_sys_tmp2214;
	wire signed [31:0] w_sys_tmp2225;
	wire signed [31:0] w_sys_tmp2226;
	wire signed [31:0] w_sys_tmp2237;
	wire signed [31:0] w_sys_tmp2238;
	wire signed [31:0] w_sys_tmp2249;
	wire signed [31:0] w_sys_tmp2250;
	wire signed [31:0] w_sys_tmp2261;
	wire signed [31:0] w_sys_tmp2262;
	wire signed [31:0] w_sys_tmp2273;
	wire signed [31:0] w_sys_tmp2274;
	wire signed [31:0] w_sys_tmp2285;
	wire signed [31:0] w_sys_tmp2286;
	wire signed [31:0] w_sys_tmp2297;
	wire signed [31:0] w_sys_tmp2298;
	wire signed [31:0] w_sys_tmp2309;
	wire signed [31:0] w_sys_tmp2310;
	wire signed [31:0] w_sys_tmp2321;
	wire signed [31:0] w_sys_tmp2322;
	wire signed [31:0] w_sys_tmp2333;
	wire signed [31:0] w_sys_tmp2334;
	wire signed [31:0] w_sys_tmp2345;
	wire signed [31:0] w_sys_tmp2346;
	wire signed [31:0] w_sys_tmp2357;
	wire signed [31:0] w_sys_tmp2358;
	wire signed [31:0] w_sys_tmp2369;
	wire signed [31:0] w_sys_tmp2370;
	wire signed [31:0] w_sys_tmp2381;
	wire signed [31:0] w_sys_tmp2382;
	wire signed [31:0] w_sys_tmp2393;
	wire signed [31:0] w_sys_tmp2394;
	wire signed [31:0] w_sys_tmp2429;
	wire signed [31:0] w_sys_tmp2430;
	wire signed [31:0] w_sys_tmp2441;
	wire signed [31:0] w_sys_tmp2442;
	wire signed [31:0] w_sys_tmp2453;
	wire signed [31:0] w_sys_tmp2454;
	wire signed [31:0] w_sys_tmp2465;
	wire signed [31:0] w_sys_tmp2466;
	wire signed [31:0] w_sys_tmp2477;
	wire signed [31:0] w_sys_tmp2478;
	wire signed [31:0] w_sys_tmp2489;
	wire signed [31:0] w_sys_tmp2490;
	wire signed [31:0] w_sys_tmp2501;
	wire signed [31:0] w_sys_tmp2502;
	wire signed [31:0] w_sys_tmp2513;
	wire signed [31:0] w_sys_tmp2514;
	wire signed [31:0] w_sys_tmp2525;
	wire signed [31:0] w_sys_tmp2526;
	wire signed [31:0] w_sys_tmp2537;
	wire signed [31:0] w_sys_tmp2538;
	wire signed [31:0] w_sys_tmp2549;
	wire signed [31:0] w_sys_tmp2550;
	wire signed [31:0] w_sys_tmp2561;
	wire signed [31:0] w_sys_tmp2562;
	wire signed [31:0] w_sys_tmp2573;
	wire signed [31:0] w_sys_tmp2574;
	wire signed [31:0] w_sys_tmp2585;
	wire signed [31:0] w_sys_tmp2586;
	wire signed [31:0] w_sys_tmp2597;
	wire signed [31:0] w_sys_tmp2598;
	wire signed [31:0] w_sys_tmp2609;
	wire signed [31:0] w_sys_tmp2610;
	wire signed [31:0] w_sys_tmp2621;
	wire signed [31:0] w_sys_tmp2622;
	wire signed [31:0] w_sys_tmp2633;
	wire signed [31:0] w_sys_tmp2634;
	wire signed [31:0] w_sys_tmp2645;
	wire signed [31:0] w_sys_tmp2646;
	wire signed [31:0] w_sys_tmp2657;
	wire signed [31:0] w_sys_tmp2658;
	wire signed [31:0] w_sys_tmp2681;
	wire signed [31:0] w_sys_tmp2682;
	wire signed [31:0] w_sys_tmp2693;
	wire signed [31:0] w_sys_tmp2694;
	wire signed [31:0] w_sys_tmp2705;
	wire signed [31:0] w_sys_tmp2706;
	wire signed [31:0] w_sys_tmp2717;
	wire signed [31:0] w_sys_tmp2718;
	wire signed [31:0] w_sys_tmp2729;
	wire signed [31:0] w_sys_tmp2730;
	wire signed [31:0] w_sys_tmp2741;
	wire signed [31:0] w_sys_tmp2742;
	wire signed [31:0] w_sys_tmp2753;
	wire signed [31:0] w_sys_tmp2754;
	wire signed [31:0] w_sys_tmp2765;
	wire signed [31:0] w_sys_tmp2766;
	wire signed [31:0] w_sys_tmp2777;
	wire signed [31:0] w_sys_tmp2778;
	wire signed [31:0] w_sys_tmp2789;
	wire signed [31:0] w_sys_tmp2790;
	wire signed [31:0] w_sys_tmp2801;
	wire signed [31:0] w_sys_tmp2802;
	wire signed [31:0] w_sys_tmp2813;
	wire signed [31:0] w_sys_tmp2814;
	wire signed [31:0] w_sys_tmp2825;
	wire signed [31:0] w_sys_tmp2826;
	wire signed [31:0] w_sys_tmp2837;
	wire signed [31:0] w_sys_tmp2838;
	wire signed [31:0] w_sys_tmp2849;
	wire signed [31:0] w_sys_tmp2850;
	wire signed [31:0] w_sys_tmp2861;
	wire signed [31:0] w_sys_tmp2862;
	wire signed [31:0] w_sys_tmp2873;
	wire signed [31:0] w_sys_tmp2874;
	wire signed [31:0] w_sys_tmp2885;
	wire signed [31:0] w_sys_tmp2886;
	wire signed [31:0] w_sys_tmp2897;
	wire signed [31:0] w_sys_tmp2898;
	wire signed [31:0] w_sys_tmp2909;
	wire signed [31:0] w_sys_tmp2910;
	wire signed [31:0] w_sys_tmp2945;
	wire signed [31:0] w_sys_tmp2946;
	wire signed [31:0] w_sys_tmp2957;
	wire signed [31:0] w_sys_tmp2958;
	wire signed [31:0] w_sys_tmp2969;
	wire signed [31:0] w_sys_tmp2970;
	wire signed [31:0] w_sys_tmp2981;
	wire signed [31:0] w_sys_tmp2982;
	wire signed [31:0] w_sys_tmp2993;
	wire signed [31:0] w_sys_tmp2994;
	wire signed [31:0] w_sys_tmp3005;
	wire signed [31:0] w_sys_tmp3006;
	wire signed [31:0] w_sys_tmp3017;
	wire signed [31:0] w_sys_tmp3018;
	wire signed [31:0] w_sys_tmp3029;
	wire signed [31:0] w_sys_tmp3030;
	wire signed [31:0] w_sys_tmp3041;
	wire signed [31:0] w_sys_tmp3042;
	wire signed [31:0] w_sys_tmp3053;
	wire signed [31:0] w_sys_tmp3054;
	wire signed [31:0] w_sys_tmp3065;
	wire signed [31:0] w_sys_tmp3066;
	wire signed [31:0] w_sys_tmp3077;
	wire signed [31:0] w_sys_tmp3078;
	wire signed [31:0] w_sys_tmp3089;
	wire signed [31:0] w_sys_tmp3090;
	wire signed [31:0] w_sys_tmp3101;
	wire signed [31:0] w_sys_tmp3102;
	wire signed [31:0] w_sys_tmp3113;
	wire signed [31:0] w_sys_tmp3114;
	wire signed [31:0] w_sys_tmp3125;
	wire signed [31:0] w_sys_tmp3126;
	wire signed [31:0] w_sys_tmp3137;
	wire signed [31:0] w_sys_tmp3138;
	wire signed [31:0] w_sys_tmp3149;
	wire signed [31:0] w_sys_tmp3150;
	wire signed [31:0] w_sys_tmp3161;
	wire signed [31:0] w_sys_tmp3162;
	wire signed [31:0] w_sys_tmp3173;
	wire signed [31:0] w_sys_tmp3174;
	wire signed [31:0] w_sys_tmp3185;
	wire signed [31:0] w_sys_tmp3186;
	wire signed [31:0] w_sys_tmp3197;
	wire signed [31:0] w_sys_tmp3198;
	wire signed [31:0] w_sys_tmp3209;
	wire signed [31:0] w_sys_tmp3210;
	wire signed [31:0] w_sys_tmp3221;
	wire signed [31:0] w_sys_tmp3222;
	wire signed [31:0] w_sys_tmp3233;
	wire signed [31:0] w_sys_tmp3234;
	wire signed [31:0] w_sys_tmp3245;
	wire signed [31:0] w_sys_tmp3246;
	wire signed [31:0] w_sys_tmp3257;
	wire signed [31:0] w_sys_tmp3258;
	wire signed [31:0] w_sys_tmp3269;
	wire signed [31:0] w_sys_tmp3270;
	wire signed [31:0] w_sys_tmp3281;
	wire signed [31:0] w_sys_tmp3282;
	wire signed [31:0] w_sys_tmp3293;
	wire signed [31:0] w_sys_tmp3294;
	wire signed [31:0] w_sys_tmp3305;
	wire signed [31:0] w_sys_tmp3306;
	wire signed [31:0] w_sys_tmp3317;
	wire signed [31:0] w_sys_tmp3318;
	wire signed [31:0] w_sys_tmp3329;
	wire signed [31:0] w_sys_tmp3330;
	wire signed [31:0] w_sys_tmp3341;
	wire signed [31:0] w_sys_tmp3342;
	wire signed [31:0] w_sys_tmp3353;
	wire signed [31:0] w_sys_tmp3354;
	wire signed [31:0] w_sys_tmp3365;
	wire signed [31:0] w_sys_tmp3366;
	wire signed [31:0] w_sys_tmp3377;
	wire signed [31:0] w_sys_tmp3378;
	wire signed [31:0] w_sys_tmp3389;
	wire signed [31:0] w_sys_tmp3390;
	wire signed [31:0] w_sys_tmp3401;
	wire signed [31:0] w_sys_tmp3402;
	wire signed [31:0] w_sys_tmp3413;
	wire signed [31:0] w_sys_tmp3414;
	wire signed [31:0] w_sys_tmp3437;
	wire signed [31:0] w_sys_tmp3438;
	wire signed [31:0] w_sys_tmp3449;
	wire signed [31:0] w_sys_tmp3450;
	wire signed [31:0] w_sys_tmp3461;
	wire signed [31:0] w_sys_tmp3462;
	wire signed [31:0] w_sys_tmp3473;
	wire signed [31:0] w_sys_tmp3474;
	wire signed [31:0] w_sys_tmp3485;
	wire signed [31:0] w_sys_tmp3486;
	wire signed [31:0] w_sys_tmp3497;
	wire signed [31:0] w_sys_tmp3498;
	wire signed [31:0] w_sys_tmp3509;
	wire signed [31:0] w_sys_tmp3510;
	wire signed [31:0] w_sys_tmp3521;
	wire signed [31:0] w_sys_tmp3522;
	wire signed [31:0] w_sys_tmp3533;
	wire signed [31:0] w_sys_tmp3534;
	wire signed [31:0] w_sys_tmp3545;
	wire signed [31:0] w_sys_tmp3546;
	wire signed [31:0] w_sys_tmp3557;
	wire signed [31:0] w_sys_tmp3558;
	wire signed [31:0] w_sys_tmp3569;
	wire signed [31:0] w_sys_tmp3570;
	wire signed [31:0] w_sys_tmp3581;
	wire signed [31:0] w_sys_tmp3582;
	wire signed [31:0] w_sys_tmp3593;
	wire signed [31:0] w_sys_tmp3594;
	wire signed [31:0] w_sys_tmp3605;
	wire signed [31:0] w_sys_tmp3606;
	wire signed [31:0] w_sys_tmp3617;
	wire signed [31:0] w_sys_tmp3618;
	wire signed [31:0] w_sys_tmp3629;
	wire signed [31:0] w_sys_tmp3630;
	wire signed [31:0] w_sys_tmp3641;
	wire signed [31:0] w_sys_tmp3642;
	wire signed [31:0] w_sys_tmp3653;
	wire signed [31:0] w_sys_tmp3654;
	wire signed [31:0] w_sys_tmp3665;
	wire signed [31:0] w_sys_tmp3666;
	wire signed [31:0] w_sys_tmp3677;
	wire signed [31:0] w_sys_tmp3678;
	wire signed [31:0] w_sys_tmp3713;
	wire signed [31:0] w_sys_tmp3714;
	wire signed [31:0] w_sys_tmp3725;
	wire signed [31:0] w_sys_tmp3726;
	wire signed [31:0] w_sys_tmp3737;
	wire signed [31:0] w_sys_tmp3738;
	wire signed [31:0] w_sys_tmp3749;
	wire signed [31:0] w_sys_tmp3750;
	wire signed [31:0] w_sys_tmp3761;
	wire signed [31:0] w_sys_tmp3762;
	wire signed [31:0] w_sys_tmp3773;
	wire signed [31:0] w_sys_tmp3774;
	wire signed [31:0] w_sys_tmp3785;
	wire signed [31:0] w_sys_tmp3786;
	wire signed [31:0] w_sys_tmp3797;
	wire signed [31:0] w_sys_tmp3798;
	wire signed [31:0] w_sys_tmp3809;
	wire signed [31:0] w_sys_tmp3810;
	wire signed [31:0] w_sys_tmp3821;
	wire signed [31:0] w_sys_tmp3822;
	wire signed [31:0] w_sys_tmp3833;
	wire signed [31:0] w_sys_tmp3834;
	wire signed [31:0] w_sys_tmp3845;
	wire signed [31:0] w_sys_tmp3846;
	wire signed [31:0] w_sys_tmp3857;
	wire signed [31:0] w_sys_tmp3858;
	wire signed [31:0] w_sys_tmp3869;
	wire signed [31:0] w_sys_tmp3870;
	wire signed [31:0] w_sys_tmp3881;
	wire signed [31:0] w_sys_tmp3882;
	wire signed [31:0] w_sys_tmp3893;
	wire signed [31:0] w_sys_tmp3894;
	wire signed [31:0] w_sys_tmp3905;
	wire signed [31:0] w_sys_tmp3906;
	wire signed [31:0] w_sys_tmp3917;
	wire signed [31:0] w_sys_tmp3918;
	wire signed [31:0] w_sys_tmp3929;
	wire signed [31:0] w_sys_tmp3930;
	wire signed [31:0] w_sys_tmp3941;
	wire signed [31:0] w_sys_tmp3942;
	wire signed [31:0] w_sys_tmp3965;
	wire signed [31:0] w_sys_tmp3966;
	wire signed [31:0] w_sys_tmp3977;
	wire signed [31:0] w_sys_tmp3978;
	wire signed [31:0] w_sys_tmp3989;
	wire signed [31:0] w_sys_tmp3990;
	wire signed [31:0] w_sys_tmp4001;
	wire signed [31:0] w_sys_tmp4002;
	wire signed [31:0] w_sys_tmp4013;
	wire signed [31:0] w_sys_tmp4014;
	wire signed [31:0] w_sys_tmp4025;
	wire signed [31:0] w_sys_tmp4026;
	wire signed [31:0] w_sys_tmp4037;
	wire signed [31:0] w_sys_tmp4038;
	wire signed [31:0] w_sys_tmp4049;
	wire signed [31:0] w_sys_tmp4050;
	wire signed [31:0] w_sys_tmp4061;
	wire signed [31:0] w_sys_tmp4062;
	wire signed [31:0] w_sys_tmp4073;
	wire signed [31:0] w_sys_tmp4074;
	wire signed [31:0] w_sys_tmp4085;
	wire signed [31:0] w_sys_tmp4086;
	wire signed [31:0] w_sys_tmp4097;
	wire signed [31:0] w_sys_tmp4098;
	wire signed [31:0] w_sys_tmp4109;
	wire signed [31:0] w_sys_tmp4110;
	wire signed [31:0] w_sys_tmp4121;
	wire signed [31:0] w_sys_tmp4122;
	wire signed [31:0] w_sys_tmp4133;
	wire signed [31:0] w_sys_tmp4134;
	wire signed [31:0] w_sys_tmp4145;
	wire signed [31:0] w_sys_tmp4146;
	wire signed [31:0] w_sys_tmp4157;
	wire signed [31:0] w_sys_tmp4158;
	wire signed [31:0] w_sys_tmp4169;
	wire signed [31:0] w_sys_tmp4170;
	wire signed [31:0] w_sys_tmp4181;
	wire signed [31:0] w_sys_tmp4182;
	wire signed [31:0] w_sys_tmp4193;
	wire signed [31:0] w_sys_tmp4194;
	wire signed [31:0] w_sys_tmp4229;
	wire signed [31:0] w_sys_tmp4230;
	wire signed [31:0] w_sys_tmp4241;
	wire signed [31:0] w_sys_tmp4242;
	wire signed [31:0] w_sys_tmp4253;
	wire signed [31:0] w_sys_tmp4254;
	wire signed [31:0] w_sys_tmp4265;
	wire signed [31:0] w_sys_tmp4266;
	wire signed [31:0] w_sys_tmp4277;
	wire signed [31:0] w_sys_tmp4278;
	wire signed [31:0] w_sys_tmp4289;
	wire signed [31:0] w_sys_tmp4290;
	wire signed [31:0] w_sys_tmp4301;
	wire signed [31:0] w_sys_tmp4302;
	wire signed [31:0] w_sys_tmp4313;
	wire signed [31:0] w_sys_tmp4314;
	wire signed [31:0] w_sys_tmp4325;
	wire signed [31:0] w_sys_tmp4326;
	wire signed [31:0] w_sys_tmp4337;
	wire signed [31:0] w_sys_tmp4338;
	wire signed [31:0] w_sys_tmp4349;
	wire signed [31:0] w_sys_tmp4350;
	wire signed [31:0] w_sys_tmp4361;
	wire signed [31:0] w_sys_tmp4362;
	wire signed [31:0] w_sys_tmp4373;
	wire signed [31:0] w_sys_tmp4374;
	wire signed [31:0] w_sys_tmp4385;
	wire signed [31:0] w_sys_tmp4386;
	wire signed [31:0] w_sys_tmp4397;
	wire signed [31:0] w_sys_tmp4398;
	wire signed [31:0] w_sys_tmp4409;
	wire signed [31:0] w_sys_tmp4410;
	wire signed [31:0] w_sys_tmp4421;
	wire signed [31:0] w_sys_tmp4422;
	wire signed [31:0] w_sys_tmp4433;
	wire signed [31:0] w_sys_tmp4434;
	wire signed [31:0] w_sys_tmp4445;
	wire signed [31:0] w_sys_tmp4446;
	wire signed [31:0] w_sys_tmp4457;
	wire signed [31:0] w_sys_tmp4458;
	wire signed [31:0] w_sys_tmp4469;
	wire signed [31:0] w_sys_tmp4470;
	wire signed [31:0] w_sys_tmp4481;
	wire signed [31:0] w_sys_tmp4482;
	wire signed [31:0] w_sys_tmp4493;
	wire signed [31:0] w_sys_tmp4494;
	wire signed [31:0] w_sys_tmp4505;
	wire signed [31:0] w_sys_tmp4506;
	wire signed [31:0] w_sys_tmp4517;
	wire signed [31:0] w_sys_tmp4518;
	wire signed [31:0] w_sys_tmp4529;
	wire signed [31:0] w_sys_tmp4530;
	wire signed [31:0] w_sys_tmp4541;
	wire signed [31:0] w_sys_tmp4542;
	wire signed [31:0] w_sys_tmp4553;
	wire signed [31:0] w_sys_tmp4554;
	wire signed [31:0] w_sys_tmp4565;
	wire signed [31:0] w_sys_tmp4566;
	wire signed [31:0] w_sys_tmp4577;
	wire signed [31:0] w_sys_tmp4578;
	wire signed [31:0] w_sys_tmp4589;
	wire signed [31:0] w_sys_tmp4590;
	wire signed [31:0] w_sys_tmp4601;
	wire signed [31:0] w_sys_tmp4602;
	wire signed [31:0] w_sys_tmp4613;
	wire signed [31:0] w_sys_tmp4614;
	wire signed [31:0] w_sys_tmp4625;
	wire signed [31:0] w_sys_tmp4626;
	wire signed [31:0] w_sys_tmp4637;
	wire signed [31:0] w_sys_tmp4638;
	wire signed [31:0] w_sys_tmp4649;
	wire signed [31:0] w_sys_tmp4650;
	wire signed [31:0] w_sys_tmp4661;
	wire signed [31:0] w_sys_tmp4662;
	wire signed [31:0] w_sys_tmp4673;
	wire signed [31:0] w_sys_tmp4674;
	wire signed [31:0] w_sys_tmp4685;
	wire signed [31:0] w_sys_tmp4686;
	wire signed [31:0] w_sys_tmp4697;
	wire signed [31:0] w_sys_tmp4698;
	wire signed [31:0] w_sys_tmp4721;
	wire signed [31:0] w_sys_tmp4722;
	wire signed [31:0] w_sys_tmp4733;
	wire signed [31:0] w_sys_tmp4734;
	wire signed [31:0] w_sys_tmp4745;
	wire signed [31:0] w_sys_tmp4746;
	wire signed [31:0] w_sys_tmp4757;
	wire signed [31:0] w_sys_tmp4758;
	wire signed [31:0] w_sys_tmp4769;
	wire signed [31:0] w_sys_tmp4770;
	wire signed [31:0] w_sys_tmp4781;
	wire signed [31:0] w_sys_tmp4782;
	wire signed [31:0] w_sys_tmp4793;
	wire signed [31:0] w_sys_tmp4794;
	wire signed [31:0] w_sys_tmp4805;
	wire signed [31:0] w_sys_tmp4806;
	wire signed [31:0] w_sys_tmp4817;
	wire signed [31:0] w_sys_tmp4818;
	wire signed [31:0] w_sys_tmp4829;
	wire signed [31:0] w_sys_tmp4830;
	wire signed [31:0] w_sys_tmp4841;
	wire signed [31:0] w_sys_tmp4842;
	wire signed [31:0] w_sys_tmp4853;
	wire signed [31:0] w_sys_tmp4854;
	wire signed [31:0] w_sys_tmp4865;
	wire signed [31:0] w_sys_tmp4866;
	wire signed [31:0] w_sys_tmp4877;
	wire signed [31:0] w_sys_tmp4878;
	wire signed [31:0] w_sys_tmp4889;
	wire signed [31:0] w_sys_tmp4890;
	wire signed [31:0] w_sys_tmp4901;
	wire signed [31:0] w_sys_tmp4902;
	wire signed [31:0] w_sys_tmp4913;
	wire signed [31:0] w_sys_tmp4914;
	wire signed [31:0] w_sys_tmp4925;
	wire signed [31:0] w_sys_tmp4926;
	wire signed [31:0] w_sys_tmp4937;
	wire signed [31:0] w_sys_tmp4938;
	wire signed [31:0] w_sys_tmp4949;
	wire signed [31:0] w_sys_tmp4950;
	wire signed [31:0] w_sys_tmp4961;
	wire signed [31:0] w_sys_tmp4962;
	wire signed [31:0] w_sys_tmp4997;
	wire signed [31:0] w_sys_tmp4998;
	wire signed [31:0] w_sys_tmp5009;
	wire signed [31:0] w_sys_tmp5010;
	wire signed [31:0] w_sys_tmp5021;
	wire signed [31:0] w_sys_tmp5022;
	wire signed [31:0] w_sys_tmp5033;
	wire signed [31:0] w_sys_tmp5034;
	wire signed [31:0] w_sys_tmp5045;
	wire signed [31:0] w_sys_tmp5046;
	wire signed [31:0] w_sys_tmp5057;
	wire signed [31:0] w_sys_tmp5058;
	wire signed [31:0] w_sys_tmp5069;
	wire signed [31:0] w_sys_tmp5070;
	wire signed [31:0] w_sys_tmp5081;
	wire signed [31:0] w_sys_tmp5082;
	wire signed [31:0] w_sys_tmp5093;
	wire signed [31:0] w_sys_tmp5094;
	wire signed [31:0] w_sys_tmp5105;
	wire signed [31:0] w_sys_tmp5106;
	wire signed [31:0] w_sys_tmp5117;
	wire signed [31:0] w_sys_tmp5118;
	wire signed [31:0] w_sys_tmp5129;
	wire signed [31:0] w_sys_tmp5130;
	wire signed [31:0] w_sys_tmp5141;
	wire signed [31:0] w_sys_tmp5142;
	wire signed [31:0] w_sys_tmp5153;
	wire signed [31:0] w_sys_tmp5154;
	wire signed [31:0] w_sys_tmp5165;
	wire signed [31:0] w_sys_tmp5166;
	wire signed [31:0] w_sys_tmp5177;
	wire signed [31:0] w_sys_tmp5178;
	wire signed [31:0] w_sys_tmp5189;
	wire signed [31:0] w_sys_tmp5190;
	wire signed [31:0] w_sys_tmp5201;
	wire signed [31:0] w_sys_tmp5202;
	wire signed [31:0] w_sys_tmp5213;
	wire signed [31:0] w_sys_tmp5214;
	wire signed [31:0] w_sys_tmp5225;
	wire signed [31:0] w_sys_tmp5226;
	wire signed [31:0] w_sys_tmp5261;
	wire signed [31:0] w_sys_tmp5262;
	wire signed [31:0] w_sys_tmp5273;
	wire signed [31:0] w_sys_tmp5274;
	wire signed [31:0] w_sys_tmp5285;
	wire signed [31:0] w_sys_tmp5286;
	wire signed [31:0] w_sys_tmp5297;
	wire signed [31:0] w_sys_tmp5298;
	wire signed [31:0] w_sys_tmp5309;
	wire signed [31:0] w_sys_tmp5310;
	wire signed [31:0] w_sys_tmp5321;
	wire signed [31:0] w_sys_tmp5322;
	wire signed [31:0] w_sys_tmp5333;
	wire signed [31:0] w_sys_tmp5334;
	wire signed [31:0] w_sys_tmp5345;
	wire signed [31:0] w_sys_tmp5346;
	wire signed [31:0] w_sys_tmp5357;
	wire signed [31:0] w_sys_tmp5358;
	wire signed [31:0] w_sys_tmp5369;
	wire signed [31:0] w_sys_tmp5370;
	wire signed [31:0] w_sys_tmp5381;
	wire signed [31:0] w_sys_tmp5382;
	wire signed [31:0] w_sys_tmp5393;
	wire signed [31:0] w_sys_tmp5394;
	wire signed [31:0] w_sys_tmp5405;
	wire signed [31:0] w_sys_tmp5406;
	wire signed [31:0] w_sys_tmp5417;
	wire signed [31:0] w_sys_tmp5418;
	wire signed [31:0] w_sys_tmp5429;
	wire signed [31:0] w_sys_tmp5430;
	wire signed [31:0] w_sys_tmp5441;
	wire signed [31:0] w_sys_tmp5442;
	wire signed [31:0] w_sys_tmp5453;
	wire signed [31:0] w_sys_tmp5454;
	wire signed [31:0] w_sys_tmp5465;
	wire signed [31:0] w_sys_tmp5466;
	wire signed [31:0] w_sys_tmp5477;
	wire signed [31:0] w_sys_tmp5478;
	wire signed [31:0] w_sys_tmp5489;
	wire signed [31:0] w_sys_tmp5490;
	wire signed [31:0] w_sys_tmp5525;
	wire signed [31:0] w_sys_tmp5526;
	wire signed [31:0] w_sys_tmp5537;
	wire signed [31:0] w_sys_tmp5538;
	wire signed [31:0] w_sys_tmp5549;
	wire signed [31:0] w_sys_tmp5550;
	wire signed [31:0] w_sys_tmp5561;
	wire signed [31:0] w_sys_tmp5562;
	wire signed [31:0] w_sys_tmp5573;
	wire signed [31:0] w_sys_tmp5574;
	wire signed [31:0] w_sys_tmp5585;
	wire signed [31:0] w_sys_tmp5586;
	wire signed [31:0] w_sys_tmp5597;
	wire signed [31:0] w_sys_tmp5598;
	wire signed [31:0] w_sys_tmp5609;
	wire signed [31:0] w_sys_tmp5610;
	wire signed [31:0] w_sys_tmp5621;
	wire signed [31:0] w_sys_tmp5622;
	wire signed [31:0] w_sys_tmp5633;
	wire signed [31:0] w_sys_tmp5634;
	wire signed [31:0] w_sys_tmp5645;
	wire signed [31:0] w_sys_tmp5646;
	wire signed [31:0] w_sys_tmp5657;
	wire signed [31:0] w_sys_tmp5658;
	wire signed [31:0] w_sys_tmp5669;
	wire signed [31:0] w_sys_tmp5670;
	wire signed [31:0] w_sys_tmp5681;
	wire signed [31:0] w_sys_tmp5682;
	wire signed [31:0] w_sys_tmp5693;
	wire signed [31:0] w_sys_tmp5694;
	wire signed [31:0] w_sys_tmp5705;
	wire signed [31:0] w_sys_tmp5706;
	wire signed [31:0] w_sys_tmp5717;
	wire signed [31:0] w_sys_tmp5718;
	wire signed [31:0] w_sys_tmp5729;
	wire signed [31:0] w_sys_tmp5730;
	wire signed [31:0] w_sys_tmp5741;
	wire signed [31:0] w_sys_tmp5742;
	wire signed [31:0] w_sys_tmp5752;
	wire signed [31:0] w_sys_tmp5753;
	wire               w_sys_tmp5754;
	wire               w_sys_tmp5755;
	wire signed [31:0] w_sys_tmp5756;
	wire signed [31:0] w_sys_tmp5759;
	wire signed [31:0] w_sys_tmp5760;
	wire        [31:0] w_sys_tmp5761;
	wire        [31:0] w_sys_tmp5767;
	wire signed [31:0] w_sys_tmp5771;
	wire signed [31:0] w_sys_tmp5772;
	wire signed [31:0] w_sys_tmp5783;
	wire signed [31:0] w_sys_tmp5784;
	wire signed [31:0] w_sys_tmp5795;
	wire signed [31:0] w_sys_tmp5796;
	wire signed [31:0] w_sys_tmp5807;
	wire signed [31:0] w_sys_tmp5808;
	wire signed [31:0] w_sys_tmp5819;
	wire signed [31:0] w_sys_tmp5820;
	wire signed [31:0] w_sys_tmp5831;
	wire signed [31:0] w_sys_tmp5832;
	wire signed [31:0] w_sys_tmp5843;
	wire signed [31:0] w_sys_tmp5844;
	wire signed [31:0] w_sys_tmp5855;
	wire signed [31:0] w_sys_tmp5856;
	wire signed [31:0] w_sys_tmp5867;
	wire signed [31:0] w_sys_tmp5868;
	wire signed [31:0] w_sys_tmp5879;
	wire signed [31:0] w_sys_tmp5880;
	wire signed [31:0] w_sys_tmp5891;
	wire signed [31:0] w_sys_tmp5892;
	wire signed [31:0] w_sys_tmp5903;
	wire signed [31:0] w_sys_tmp5904;
	wire signed [31:0] w_sys_tmp5915;
	wire signed [31:0] w_sys_tmp5916;
	wire signed [31:0] w_sys_tmp5927;
	wire signed [31:0] w_sys_tmp5928;
	wire signed [31:0] w_sys_tmp5939;
	wire signed [31:0] w_sys_tmp5940;
	wire signed [31:0] w_sys_tmp5951;
	wire signed [31:0] w_sys_tmp5952;
	wire signed [31:0] w_sys_tmp5963;
	wire signed [31:0] w_sys_tmp5964;
	wire signed [31:0] w_sys_tmp5975;
	wire signed [31:0] w_sys_tmp5976;
	wire signed [31:0] w_sys_tmp5987;
	wire signed [31:0] w_sys_tmp5988;
	wire signed [31:0] w_sys_tmp5999;
	wire signed [31:0] w_sys_tmp6000;
	wire signed [31:0] w_sys_tmp6023;
	wire signed [31:0] w_sys_tmp6024;
	wire signed [31:0] w_sys_tmp6035;
	wire signed [31:0] w_sys_tmp6036;
	wire signed [31:0] w_sys_tmp6047;
	wire signed [31:0] w_sys_tmp6048;
	wire signed [31:0] w_sys_tmp6059;
	wire signed [31:0] w_sys_tmp6060;
	wire signed [31:0] w_sys_tmp6071;
	wire signed [31:0] w_sys_tmp6072;
	wire signed [31:0] w_sys_tmp6083;
	wire signed [31:0] w_sys_tmp6084;
	wire signed [31:0] w_sys_tmp6095;
	wire signed [31:0] w_sys_tmp6096;
	wire signed [31:0] w_sys_tmp6107;
	wire signed [31:0] w_sys_tmp6108;
	wire signed [31:0] w_sys_tmp6119;
	wire signed [31:0] w_sys_tmp6120;
	wire signed [31:0] w_sys_tmp6131;
	wire signed [31:0] w_sys_tmp6132;
	wire signed [31:0] w_sys_tmp6143;
	wire signed [31:0] w_sys_tmp6144;
	wire signed [31:0] w_sys_tmp6155;
	wire signed [31:0] w_sys_tmp6156;
	wire signed [31:0] w_sys_tmp6167;
	wire signed [31:0] w_sys_tmp6168;
	wire signed [31:0] w_sys_tmp6179;
	wire signed [31:0] w_sys_tmp6180;
	wire signed [31:0] w_sys_tmp6191;
	wire signed [31:0] w_sys_tmp6192;
	wire signed [31:0] w_sys_tmp6203;
	wire signed [31:0] w_sys_tmp6204;
	wire signed [31:0] w_sys_tmp6215;
	wire signed [31:0] w_sys_tmp6216;
	wire signed [31:0] w_sys_tmp6227;
	wire signed [31:0] w_sys_tmp6228;
	wire signed [31:0] w_sys_tmp6239;
	wire signed [31:0] w_sys_tmp6240;
	wire signed [31:0] w_sys_tmp6251;
	wire signed [31:0] w_sys_tmp6252;
	wire signed [31:0] w_sys_tmp6263;
	wire signed [31:0] w_sys_tmp6264;
	wire signed [31:0] w_sys_tmp6299;
	wire signed [31:0] w_sys_tmp6300;
	wire signed [31:0] w_sys_tmp6311;
	wire signed [31:0] w_sys_tmp6312;
	wire signed [31:0] w_sys_tmp6323;
	wire signed [31:0] w_sys_tmp6324;
	wire signed [31:0] w_sys_tmp6335;
	wire signed [31:0] w_sys_tmp6336;
	wire signed [31:0] w_sys_tmp6347;
	wire signed [31:0] w_sys_tmp6348;
	wire signed [31:0] w_sys_tmp6359;
	wire signed [31:0] w_sys_tmp6360;
	wire signed [31:0] w_sys_tmp6371;
	wire signed [31:0] w_sys_tmp6372;
	wire signed [31:0] w_sys_tmp6383;
	wire signed [31:0] w_sys_tmp6384;
	wire signed [31:0] w_sys_tmp6395;
	wire signed [31:0] w_sys_tmp6396;
	wire signed [31:0] w_sys_tmp6407;
	wire signed [31:0] w_sys_tmp6408;
	wire signed [31:0] w_sys_tmp6419;
	wire signed [31:0] w_sys_tmp6420;
	wire signed [31:0] w_sys_tmp6431;
	wire signed [31:0] w_sys_tmp6432;
	wire signed [31:0] w_sys_tmp6443;
	wire signed [31:0] w_sys_tmp6444;
	wire signed [31:0] w_sys_tmp6455;
	wire signed [31:0] w_sys_tmp6456;
	wire signed [31:0] w_sys_tmp6467;
	wire signed [31:0] w_sys_tmp6468;
	wire signed [31:0] w_sys_tmp6479;
	wire signed [31:0] w_sys_tmp6480;
	wire signed [31:0] w_sys_tmp6491;
	wire signed [31:0] w_sys_tmp6492;
	wire signed [31:0] w_sys_tmp6503;
	wire signed [31:0] w_sys_tmp6504;
	wire signed [31:0] w_sys_tmp6515;
	wire signed [31:0] w_sys_tmp6516;
	wire signed [31:0] w_sys_tmp6527;
	wire signed [31:0] w_sys_tmp6528;
	wire signed [31:0] w_sys_tmp6563;
	wire signed [31:0] w_sys_tmp6564;
	wire signed [31:0] w_sys_tmp6575;
	wire signed [31:0] w_sys_tmp6576;
	wire signed [31:0] w_sys_tmp6587;
	wire signed [31:0] w_sys_tmp6588;
	wire signed [31:0] w_sys_tmp6599;
	wire signed [31:0] w_sys_tmp6600;
	wire signed [31:0] w_sys_tmp6611;
	wire signed [31:0] w_sys_tmp6612;
	wire signed [31:0] w_sys_tmp6623;
	wire signed [31:0] w_sys_tmp6624;
	wire signed [31:0] w_sys_tmp6635;
	wire signed [31:0] w_sys_tmp6636;
	wire signed [31:0] w_sys_tmp6647;
	wire signed [31:0] w_sys_tmp6648;
	wire signed [31:0] w_sys_tmp6659;
	wire signed [31:0] w_sys_tmp6660;
	wire signed [31:0] w_sys_tmp6671;
	wire signed [31:0] w_sys_tmp6672;
	wire signed [31:0] w_sys_tmp6683;
	wire signed [31:0] w_sys_tmp6684;
	wire signed [31:0] w_sys_tmp6695;
	wire signed [31:0] w_sys_tmp6696;
	wire signed [31:0] w_sys_tmp6707;
	wire signed [31:0] w_sys_tmp6708;
	wire signed [31:0] w_sys_tmp6719;
	wire signed [31:0] w_sys_tmp6720;
	wire signed [31:0] w_sys_tmp6731;
	wire signed [31:0] w_sys_tmp6732;
	wire signed [31:0] w_sys_tmp6743;
	wire signed [31:0] w_sys_tmp6744;
	wire signed [31:0] w_sys_tmp6755;
	wire signed [31:0] w_sys_tmp6756;
	wire signed [31:0] w_sys_tmp6767;
	wire signed [31:0] w_sys_tmp6768;
	wire signed [31:0] w_sys_tmp6779;
	wire signed [31:0] w_sys_tmp6780;
	wire signed [31:0] w_sys_tmp6791;
	wire signed [31:0] w_sys_tmp6792;
	wire signed [31:0] w_sys_tmp6827;
	wire signed [31:0] w_sys_tmp6828;
	wire signed [31:0] w_sys_tmp6839;
	wire signed [31:0] w_sys_tmp6840;
	wire signed [31:0] w_sys_tmp6851;
	wire signed [31:0] w_sys_tmp6852;
	wire signed [31:0] w_sys_tmp6863;
	wire signed [31:0] w_sys_tmp6864;
	wire signed [31:0] w_sys_tmp6875;
	wire signed [31:0] w_sys_tmp6876;
	wire signed [31:0] w_sys_tmp6887;
	wire signed [31:0] w_sys_tmp6888;
	wire signed [31:0] w_sys_tmp6899;
	wire signed [31:0] w_sys_tmp6900;
	wire signed [31:0] w_sys_tmp6911;
	wire signed [31:0] w_sys_tmp6912;
	wire signed [31:0] w_sys_tmp6923;
	wire signed [31:0] w_sys_tmp6924;
	wire signed [31:0] w_sys_tmp6935;
	wire signed [31:0] w_sys_tmp6936;
	wire signed [31:0] w_sys_tmp6947;
	wire signed [31:0] w_sys_tmp6948;
	wire signed [31:0] w_sys_tmp6959;
	wire signed [31:0] w_sys_tmp6960;
	wire signed [31:0] w_sys_tmp6971;
	wire signed [31:0] w_sys_tmp6972;
	wire signed [31:0] w_sys_tmp6983;
	wire signed [31:0] w_sys_tmp6984;
	wire signed [31:0] w_sys_tmp6995;
	wire signed [31:0] w_sys_tmp6996;
	wire signed [31:0] w_sys_tmp7007;
	wire signed [31:0] w_sys_tmp7008;
	wire signed [31:0] w_sys_tmp7019;
	wire signed [31:0] w_sys_tmp7020;
	wire signed [31:0] w_sys_tmp7031;
	wire signed [31:0] w_sys_tmp7032;
	wire signed [31:0] w_sys_tmp7043;
	wire signed [31:0] w_sys_tmp7044;
	wire signed [31:0] w_sys_tmp7054;
	wire               w_sys_tmp7055;
	wire               w_sys_tmp7056;
	wire signed [31:0] w_sys_tmp7057;
	wire               w_sys_tmp7058;
	wire               w_sys_tmp7059;
	wire signed [31:0] w_sys_tmp7062;
	wire signed [31:0] w_sys_tmp7063;
	wire        [31:0] w_sys_tmp7064;
	wire signed [31:0] w_sys_tmp7066;
	wire signed [31:0] w_sys_tmp7067;
	wire        [31:0] w_sys_tmp7069;
	wire signed [31:0] w_sys_tmp7070;
	wire signed [31:0] w_sys_tmp7071;
	wire signed [31:0] w_sys_tmp7072;
	wire signed [31:0] w_sys_tmp7074;
	wire               w_sys_tmp7075;
	wire               w_sys_tmp7076;
	wire signed [31:0] w_sys_tmp7079;
	wire signed [31:0] w_sys_tmp7080;
	wire signed [31:0] w_sys_tmp7081;
	wire        [31:0] w_sys_tmp7082;
	wire signed [31:0] w_sys_tmp7084;
	wire signed [31:0] w_sys_tmp7085;
	wire signed [31:0] w_sys_tmp7088;
	wire signed [31:0] w_sys_tmp7089;
	wire signed [31:0] w_sys_tmp7318;
	wire signed [31:0] w_sys_tmp7319;
	wire               w_sys_tmp7320;
	wire               w_sys_tmp7321;
	wire signed [31:0] w_sys_tmp7322;
	wire signed [31:0] w_sys_tmp7323;
	wire signed [31:0] w_sys_tmp7326;
	wire signed [31:0] w_sys_tmp7327;
	wire signed [31:0] w_sys_tmp7328;
	wire        [31:0] w_sys_tmp7329;
	wire signed [31:0] w_sys_tmp7330;
	wire               w_sys_tmp7445;
	wire               w_sys_tmp7446;
	wire signed [31:0] w_sys_tmp7447;
	wire signed [31:0] w_sys_tmp7450;
	wire signed [31:0] w_sys_tmp7451;
	wire        [31:0] w_sys_tmp7452;
	wire signed [31:0] w_sys_tmp7456;
	wire signed [31:0] w_sys_tmp7457;
	wire signed [31:0] w_sys_tmp7462;
	wire signed [31:0] w_sys_tmp7463;
	wire signed [31:0] w_sys_tmp7468;
	wire signed [31:0] w_sys_tmp7469;
	wire signed [31:0] w_sys_tmp7474;
	wire signed [31:0] w_sys_tmp7475;
	wire signed [31:0] w_sys_tmp7480;
	wire signed [31:0] w_sys_tmp7481;
	wire signed [31:0] w_sys_tmp7486;
	wire signed [31:0] w_sys_tmp7487;
	wire signed [31:0] w_sys_tmp7492;
	wire signed [31:0] w_sys_tmp7493;
	wire signed [31:0] w_sys_tmp7498;
	wire signed [31:0] w_sys_tmp7499;
	wire signed [31:0] w_sys_tmp7504;
	wire signed [31:0] w_sys_tmp7505;
	wire signed [31:0] w_sys_tmp7510;
	wire signed [31:0] w_sys_tmp7511;
	wire signed [31:0] w_sys_tmp7516;
	wire signed [31:0] w_sys_tmp7517;
	wire signed [31:0] w_sys_tmp7522;
	wire signed [31:0] w_sys_tmp7523;
	wire signed [31:0] w_sys_tmp7528;
	wire signed [31:0] w_sys_tmp7529;
	wire signed [31:0] w_sys_tmp7534;
	wire signed [31:0] w_sys_tmp7535;
	wire signed [31:0] w_sys_tmp7540;
	wire signed [31:0] w_sys_tmp7541;
	wire signed [31:0] w_sys_tmp7546;
	wire signed [31:0] w_sys_tmp7547;
	wire signed [31:0] w_sys_tmp7552;
	wire signed [31:0] w_sys_tmp7553;
	wire signed [31:0] w_sys_tmp7558;
	wire signed [31:0] w_sys_tmp7559;
	wire signed [31:0] w_sys_tmp7564;
	wire signed [31:0] w_sys_tmp7565;
	wire signed [31:0] w_sys_tmp7570;
	wire signed [31:0] w_sys_tmp7571;
	wire signed [31:0] w_sys_tmp7576;
	wire signed [31:0] w_sys_tmp7577;
	wire signed [31:0] w_sys_tmp7594;
	wire signed [31:0] w_sys_tmp7595;
	wire signed [31:0] w_sys_tmp7600;
	wire signed [31:0] w_sys_tmp7601;
	wire signed [31:0] w_sys_tmp7606;
	wire signed [31:0] w_sys_tmp7607;
	wire signed [31:0] w_sys_tmp7612;
	wire signed [31:0] w_sys_tmp7613;
	wire signed [31:0] w_sys_tmp7618;
	wire signed [31:0] w_sys_tmp7619;
	wire signed [31:0] w_sys_tmp7624;
	wire signed [31:0] w_sys_tmp7625;
	wire signed [31:0] w_sys_tmp7630;
	wire signed [31:0] w_sys_tmp7631;
	wire signed [31:0] w_sys_tmp7636;
	wire signed [31:0] w_sys_tmp7637;
	wire signed [31:0] w_sys_tmp7642;
	wire signed [31:0] w_sys_tmp7643;
	wire signed [31:0] w_sys_tmp7648;
	wire signed [31:0] w_sys_tmp7649;
	wire signed [31:0] w_sys_tmp7654;
	wire signed [31:0] w_sys_tmp7655;
	wire signed [31:0] w_sys_tmp7660;
	wire signed [31:0] w_sys_tmp7661;
	wire signed [31:0] w_sys_tmp7666;
	wire signed [31:0] w_sys_tmp7667;
	wire signed [31:0] w_sys_tmp7672;
	wire signed [31:0] w_sys_tmp7673;
	wire signed [31:0] w_sys_tmp7678;
	wire signed [31:0] w_sys_tmp7679;
	wire signed [31:0] w_sys_tmp7684;
	wire signed [31:0] w_sys_tmp7685;
	wire signed [31:0] w_sys_tmp7690;
	wire signed [31:0] w_sys_tmp7691;
	wire signed [31:0] w_sys_tmp7696;
	wire signed [31:0] w_sys_tmp7697;
	wire signed [31:0] w_sys_tmp7702;
	wire signed [31:0] w_sys_tmp7703;
	wire signed [31:0] w_sys_tmp7708;
	wire signed [31:0] w_sys_tmp7709;
	wire signed [31:0] w_sys_tmp7726;
	wire signed [31:0] w_sys_tmp7727;
	wire signed [31:0] w_sys_tmp7732;
	wire signed [31:0] w_sys_tmp7733;
	wire signed [31:0] w_sys_tmp7738;
	wire signed [31:0] w_sys_tmp7739;
	wire signed [31:0] w_sys_tmp7744;
	wire signed [31:0] w_sys_tmp7745;
	wire signed [31:0] w_sys_tmp7750;
	wire signed [31:0] w_sys_tmp7751;
	wire signed [31:0] w_sys_tmp7756;
	wire signed [31:0] w_sys_tmp7757;
	wire signed [31:0] w_sys_tmp7762;
	wire signed [31:0] w_sys_tmp7763;
	wire signed [31:0] w_sys_tmp7768;
	wire signed [31:0] w_sys_tmp7769;
	wire signed [31:0] w_sys_tmp7774;
	wire signed [31:0] w_sys_tmp7775;
	wire signed [31:0] w_sys_tmp7780;
	wire signed [31:0] w_sys_tmp7781;
	wire signed [31:0] w_sys_tmp7786;
	wire signed [31:0] w_sys_tmp7787;
	wire signed [31:0] w_sys_tmp7792;
	wire signed [31:0] w_sys_tmp7793;
	wire signed [31:0] w_sys_tmp7798;
	wire signed [31:0] w_sys_tmp7799;
	wire signed [31:0] w_sys_tmp7804;
	wire signed [31:0] w_sys_tmp7805;
	wire signed [31:0] w_sys_tmp7810;
	wire signed [31:0] w_sys_tmp7811;
	wire signed [31:0] w_sys_tmp7816;
	wire signed [31:0] w_sys_tmp7817;
	wire signed [31:0] w_sys_tmp7822;
	wire signed [31:0] w_sys_tmp7823;
	wire signed [31:0] w_sys_tmp7828;
	wire signed [31:0] w_sys_tmp7829;
	wire signed [31:0] w_sys_tmp7834;
	wire signed [31:0] w_sys_tmp7835;
	wire signed [31:0] w_sys_tmp7840;
	wire signed [31:0] w_sys_tmp7841;
	wire signed [31:0] w_sys_tmp7858;
	wire signed [31:0] w_sys_tmp7859;
	wire signed [31:0] w_sys_tmp7864;
	wire signed [31:0] w_sys_tmp7865;
	wire signed [31:0] w_sys_tmp7870;
	wire signed [31:0] w_sys_tmp7871;
	wire signed [31:0] w_sys_tmp7876;
	wire signed [31:0] w_sys_tmp7877;
	wire signed [31:0] w_sys_tmp7882;
	wire signed [31:0] w_sys_tmp7883;
	wire signed [31:0] w_sys_tmp7888;
	wire signed [31:0] w_sys_tmp7889;
	wire signed [31:0] w_sys_tmp7894;
	wire signed [31:0] w_sys_tmp7895;
	wire signed [31:0] w_sys_tmp7900;
	wire signed [31:0] w_sys_tmp7901;
	wire signed [31:0] w_sys_tmp7906;
	wire signed [31:0] w_sys_tmp7907;
	wire signed [31:0] w_sys_tmp7912;
	wire signed [31:0] w_sys_tmp7913;
	wire signed [31:0] w_sys_tmp7918;
	wire signed [31:0] w_sys_tmp7919;
	wire signed [31:0] w_sys_tmp7924;
	wire signed [31:0] w_sys_tmp7925;
	wire signed [31:0] w_sys_tmp7930;
	wire signed [31:0] w_sys_tmp7931;
	wire signed [31:0] w_sys_tmp7936;
	wire signed [31:0] w_sys_tmp7937;
	wire signed [31:0] w_sys_tmp7942;
	wire signed [31:0] w_sys_tmp7943;
	wire signed [31:0] w_sys_tmp7948;
	wire signed [31:0] w_sys_tmp7949;
	wire signed [31:0] w_sys_tmp7954;
	wire signed [31:0] w_sys_tmp7955;
	wire signed [31:0] w_sys_tmp7960;
	wire signed [31:0] w_sys_tmp7961;
	wire signed [31:0] w_sys_tmp7966;
	wire signed [31:0] w_sys_tmp7967;
	wire signed [31:0] w_sys_tmp7972;
	wire signed [31:0] w_sys_tmp7973;
	wire signed [31:0] w_sys_tmp7990;
	wire signed [31:0] w_sys_tmp7991;
	wire signed [31:0] w_sys_tmp7996;
	wire signed [31:0] w_sys_tmp7997;
	wire signed [31:0] w_sys_tmp8002;
	wire signed [31:0] w_sys_tmp8003;
	wire signed [31:0] w_sys_tmp8008;
	wire signed [31:0] w_sys_tmp8009;
	wire signed [31:0] w_sys_tmp8014;
	wire signed [31:0] w_sys_tmp8015;
	wire signed [31:0] w_sys_tmp8020;
	wire signed [31:0] w_sys_tmp8021;
	wire signed [31:0] w_sys_tmp8026;
	wire signed [31:0] w_sys_tmp8027;
	wire signed [31:0] w_sys_tmp8032;
	wire signed [31:0] w_sys_tmp8033;
	wire signed [31:0] w_sys_tmp8038;
	wire signed [31:0] w_sys_tmp8039;
	wire signed [31:0] w_sys_tmp8044;
	wire signed [31:0] w_sys_tmp8045;
	wire signed [31:0] w_sys_tmp8050;
	wire signed [31:0] w_sys_tmp8051;
	wire signed [31:0] w_sys_tmp8056;
	wire signed [31:0] w_sys_tmp8057;
	wire signed [31:0] w_sys_tmp8062;
	wire signed [31:0] w_sys_tmp8063;
	wire signed [31:0] w_sys_tmp8068;
	wire signed [31:0] w_sys_tmp8069;
	wire signed [31:0] w_sys_tmp8074;
	wire signed [31:0] w_sys_tmp8075;
	wire signed [31:0] w_sys_tmp8080;
	wire signed [31:0] w_sys_tmp8081;
	wire signed [31:0] w_sys_tmp8086;
	wire signed [31:0] w_sys_tmp8087;
	wire signed [31:0] w_sys_tmp8092;
	wire signed [31:0] w_sys_tmp8093;
	wire signed [31:0] w_sys_tmp8098;
	wire signed [31:0] w_sys_tmp8099;
	wire signed [31:0] w_sys_tmp8104;
	wire signed [31:0] w_sys_tmp8105;
	wire signed [31:0] w_sys_tmp8110;
	wire signed [31:0] w_sys_tmp8111;
	wire signed [31:0] w_sys_tmp8116;
	wire signed [31:0] w_sys_tmp8117;
	wire signed [31:0] w_sys_tmp8122;
	wire signed [31:0] w_sys_tmp8123;
	wire signed [31:0] w_sys_tmp8128;
	wire signed [31:0] w_sys_tmp8129;
	wire signed [31:0] w_sys_tmp8134;
	wire signed [31:0] w_sys_tmp8135;
	wire signed [31:0] w_sys_tmp8140;
	wire signed [31:0] w_sys_tmp8141;
	wire signed [31:0] w_sys_tmp8146;
	wire signed [31:0] w_sys_tmp8147;
	wire signed [31:0] w_sys_tmp8152;
	wire signed [31:0] w_sys_tmp8153;
	wire signed [31:0] w_sys_tmp8158;
	wire signed [31:0] w_sys_tmp8159;
	wire signed [31:0] w_sys_tmp8164;
	wire signed [31:0] w_sys_tmp8165;
	wire signed [31:0] w_sys_tmp8170;
	wire signed [31:0] w_sys_tmp8171;
	wire signed [31:0] w_sys_tmp8176;
	wire signed [31:0] w_sys_tmp8177;
	wire signed [31:0] w_sys_tmp8182;
	wire signed [31:0] w_sys_tmp8183;
	wire signed [31:0] w_sys_tmp8188;
	wire signed [31:0] w_sys_tmp8189;
	wire signed [31:0] w_sys_tmp8194;
	wire signed [31:0] w_sys_tmp8195;
	wire signed [31:0] w_sys_tmp8200;
	wire signed [31:0] w_sys_tmp8201;
	wire signed [31:0] w_sys_tmp8206;
	wire signed [31:0] w_sys_tmp8207;
	wire signed [31:0] w_sys_tmp8212;
	wire signed [31:0] w_sys_tmp8213;
	wire signed [31:0] w_sys_tmp8218;
	wire signed [31:0] w_sys_tmp8219;
	wire signed [31:0] w_sys_tmp8224;
	wire signed [31:0] w_sys_tmp8225;
	wire signed [31:0] w_sys_tmp8230;
	wire signed [31:0] w_sys_tmp8231;
	wire signed [31:0] w_sys_tmp8248;
	wire signed [31:0] w_sys_tmp8249;
	wire signed [31:0] w_sys_tmp8254;
	wire signed [31:0] w_sys_tmp8255;
	wire signed [31:0] w_sys_tmp8260;
	wire signed [31:0] w_sys_tmp8261;
	wire signed [31:0] w_sys_tmp8266;
	wire signed [31:0] w_sys_tmp8267;
	wire signed [31:0] w_sys_tmp8272;
	wire signed [31:0] w_sys_tmp8273;
	wire signed [31:0] w_sys_tmp8278;
	wire signed [31:0] w_sys_tmp8279;
	wire signed [31:0] w_sys_tmp8284;
	wire signed [31:0] w_sys_tmp8285;
	wire signed [31:0] w_sys_tmp8290;
	wire signed [31:0] w_sys_tmp8291;
	wire signed [31:0] w_sys_tmp8296;
	wire signed [31:0] w_sys_tmp8297;
	wire signed [31:0] w_sys_tmp8302;
	wire signed [31:0] w_sys_tmp8303;
	wire signed [31:0] w_sys_tmp8308;
	wire signed [31:0] w_sys_tmp8309;
	wire signed [31:0] w_sys_tmp8314;
	wire signed [31:0] w_sys_tmp8315;
	wire signed [31:0] w_sys_tmp8320;
	wire signed [31:0] w_sys_tmp8321;
	wire signed [31:0] w_sys_tmp8326;
	wire signed [31:0] w_sys_tmp8327;
	wire signed [31:0] w_sys_tmp8332;
	wire signed [31:0] w_sys_tmp8333;
	wire signed [31:0] w_sys_tmp8338;
	wire signed [31:0] w_sys_tmp8339;
	wire signed [31:0] w_sys_tmp8344;
	wire signed [31:0] w_sys_tmp8345;
	wire signed [31:0] w_sys_tmp8350;
	wire signed [31:0] w_sys_tmp8351;
	wire signed [31:0] w_sys_tmp8356;
	wire signed [31:0] w_sys_tmp8357;
	wire signed [31:0] w_sys_tmp8362;
	wire signed [31:0] w_sys_tmp8363;
	wire signed [31:0] w_sys_tmp8380;
	wire signed [31:0] w_sys_tmp8381;
	wire signed [31:0] w_sys_tmp8386;
	wire signed [31:0] w_sys_tmp8387;
	wire signed [31:0] w_sys_tmp8392;
	wire signed [31:0] w_sys_tmp8393;
	wire signed [31:0] w_sys_tmp8398;
	wire signed [31:0] w_sys_tmp8399;
	wire signed [31:0] w_sys_tmp8404;
	wire signed [31:0] w_sys_tmp8405;
	wire signed [31:0] w_sys_tmp8410;
	wire signed [31:0] w_sys_tmp8411;
	wire signed [31:0] w_sys_tmp8416;
	wire signed [31:0] w_sys_tmp8417;
	wire signed [31:0] w_sys_tmp8422;
	wire signed [31:0] w_sys_tmp8423;
	wire signed [31:0] w_sys_tmp8428;
	wire signed [31:0] w_sys_tmp8429;
	wire signed [31:0] w_sys_tmp8434;
	wire signed [31:0] w_sys_tmp8435;
	wire signed [31:0] w_sys_tmp8440;
	wire signed [31:0] w_sys_tmp8441;
	wire signed [31:0] w_sys_tmp8446;
	wire signed [31:0] w_sys_tmp8447;
	wire signed [31:0] w_sys_tmp8452;
	wire signed [31:0] w_sys_tmp8453;
	wire signed [31:0] w_sys_tmp8458;
	wire signed [31:0] w_sys_tmp8459;
	wire signed [31:0] w_sys_tmp8464;
	wire signed [31:0] w_sys_tmp8465;
	wire signed [31:0] w_sys_tmp8470;
	wire signed [31:0] w_sys_tmp8471;
	wire signed [31:0] w_sys_tmp8476;
	wire signed [31:0] w_sys_tmp8477;
	wire signed [31:0] w_sys_tmp8482;
	wire signed [31:0] w_sys_tmp8483;
	wire signed [31:0] w_sys_tmp8488;
	wire signed [31:0] w_sys_tmp8489;
	wire signed [31:0] w_sys_tmp8494;
	wire signed [31:0] w_sys_tmp8495;
	wire signed [31:0] w_sys_tmp8512;
	wire signed [31:0] w_sys_tmp8513;
	wire signed [31:0] w_sys_tmp8518;
	wire signed [31:0] w_sys_tmp8519;
	wire signed [31:0] w_sys_tmp8524;
	wire signed [31:0] w_sys_tmp8525;
	wire signed [31:0] w_sys_tmp8530;
	wire signed [31:0] w_sys_tmp8531;
	wire signed [31:0] w_sys_tmp8536;
	wire signed [31:0] w_sys_tmp8537;
	wire signed [31:0] w_sys_tmp8542;
	wire signed [31:0] w_sys_tmp8543;
	wire signed [31:0] w_sys_tmp8548;
	wire signed [31:0] w_sys_tmp8549;
	wire signed [31:0] w_sys_tmp8554;
	wire signed [31:0] w_sys_tmp8555;
	wire signed [31:0] w_sys_tmp8560;
	wire signed [31:0] w_sys_tmp8561;
	wire signed [31:0] w_sys_tmp8566;
	wire signed [31:0] w_sys_tmp8567;
	wire signed [31:0] w_sys_tmp8572;
	wire signed [31:0] w_sys_tmp8573;
	wire signed [31:0] w_sys_tmp8578;
	wire signed [31:0] w_sys_tmp8579;
	wire signed [31:0] w_sys_tmp8584;
	wire signed [31:0] w_sys_tmp8585;
	wire signed [31:0] w_sys_tmp8590;
	wire signed [31:0] w_sys_tmp8591;
	wire signed [31:0] w_sys_tmp8596;
	wire signed [31:0] w_sys_tmp8597;
	wire signed [31:0] w_sys_tmp8602;
	wire signed [31:0] w_sys_tmp8603;
	wire signed [31:0] w_sys_tmp8608;
	wire signed [31:0] w_sys_tmp8609;
	wire signed [31:0] w_sys_tmp8614;
	wire signed [31:0] w_sys_tmp8615;
	wire signed [31:0] w_sys_tmp8620;
	wire signed [31:0] w_sys_tmp8621;
	wire signed [31:0] w_sys_tmp8626;
	wire signed [31:0] w_sys_tmp8627;
	wire signed [31:0] w_sys_tmp8644;
	wire signed [31:0] w_sys_tmp8645;
	wire signed [31:0] w_sys_tmp8650;
	wire signed [31:0] w_sys_tmp8651;
	wire signed [31:0] w_sys_tmp8656;
	wire signed [31:0] w_sys_tmp8657;
	wire signed [31:0] w_sys_tmp8662;
	wire signed [31:0] w_sys_tmp8663;
	wire signed [31:0] w_sys_tmp8668;
	wire signed [31:0] w_sys_tmp8669;
	wire signed [31:0] w_sys_tmp8674;
	wire signed [31:0] w_sys_tmp8675;
	wire signed [31:0] w_sys_tmp8680;
	wire signed [31:0] w_sys_tmp8681;
	wire signed [31:0] w_sys_tmp8686;
	wire signed [31:0] w_sys_tmp8687;
	wire signed [31:0] w_sys_tmp8692;
	wire signed [31:0] w_sys_tmp8693;
	wire signed [31:0] w_sys_tmp8698;
	wire signed [31:0] w_sys_tmp8699;
	wire signed [31:0] w_sys_tmp8704;
	wire signed [31:0] w_sys_tmp8705;
	wire signed [31:0] w_sys_tmp8710;
	wire signed [31:0] w_sys_tmp8711;
	wire signed [31:0] w_sys_tmp8716;
	wire signed [31:0] w_sys_tmp8717;
	wire signed [31:0] w_sys_tmp8722;
	wire signed [31:0] w_sys_tmp8723;
	wire signed [31:0] w_sys_tmp8728;
	wire signed [31:0] w_sys_tmp8729;
	wire signed [31:0] w_sys_tmp8734;
	wire signed [31:0] w_sys_tmp8735;
	wire signed [31:0] w_sys_tmp8740;
	wire signed [31:0] w_sys_tmp8741;
	wire signed [31:0] w_sys_tmp8746;
	wire signed [31:0] w_sys_tmp8747;
	wire signed [31:0] w_sys_tmp8752;
	wire signed [31:0] w_sys_tmp8753;
	wire signed [31:0] w_sys_tmp8758;
	wire signed [31:0] w_sys_tmp8759;
	wire signed [31:0] w_sys_tmp8764;
	wire signed [31:0] w_sys_tmp8765;
	wire signed [31:0] w_sys_tmp8770;
	wire signed [31:0] w_sys_tmp8771;
	wire signed [31:0] w_sys_tmp8776;
	wire signed [31:0] w_sys_tmp8777;
	wire signed [31:0] w_sys_tmp8782;
	wire signed [31:0] w_sys_tmp8783;
	wire signed [31:0] w_sys_tmp8788;
	wire signed [31:0] w_sys_tmp8789;
	wire signed [31:0] w_sys_tmp8794;
	wire signed [31:0] w_sys_tmp8795;
	wire signed [31:0] w_sys_tmp8800;
	wire signed [31:0] w_sys_tmp8801;
	wire signed [31:0] w_sys_tmp8806;
	wire signed [31:0] w_sys_tmp8807;
	wire signed [31:0] w_sys_tmp8812;
	wire signed [31:0] w_sys_tmp8813;
	wire signed [31:0] w_sys_tmp8818;
	wire signed [31:0] w_sys_tmp8819;
	wire signed [31:0] w_sys_tmp8824;
	wire signed [31:0] w_sys_tmp8825;
	wire signed [31:0] w_sys_tmp8830;
	wire signed [31:0] w_sys_tmp8831;
	wire signed [31:0] w_sys_tmp8836;
	wire signed [31:0] w_sys_tmp8837;
	wire signed [31:0] w_sys_tmp8842;
	wire signed [31:0] w_sys_tmp8843;
	wire signed [31:0] w_sys_tmp8848;
	wire signed [31:0] w_sys_tmp8849;
	wire signed [31:0] w_sys_tmp8854;
	wire signed [31:0] w_sys_tmp8855;
	wire signed [31:0] w_sys_tmp8860;
	wire signed [31:0] w_sys_tmp8861;
	wire signed [31:0] w_sys_tmp8866;
	wire signed [31:0] w_sys_tmp8867;
	wire signed [31:0] w_sys_tmp8872;
	wire signed [31:0] w_sys_tmp8873;
	wire signed [31:0] w_sys_tmp8878;
	wire signed [31:0] w_sys_tmp8879;
	wire signed [31:0] w_sys_tmp8884;
	wire signed [31:0] w_sys_tmp8885;
	wire signed [31:0] w_sys_tmp8902;
	wire signed [31:0] w_sys_tmp8903;
	wire signed [31:0] w_sys_tmp8908;
	wire signed [31:0] w_sys_tmp8909;
	wire signed [31:0] w_sys_tmp8914;
	wire signed [31:0] w_sys_tmp8915;
	wire signed [31:0] w_sys_tmp8920;
	wire signed [31:0] w_sys_tmp8921;
	wire signed [31:0] w_sys_tmp8926;
	wire signed [31:0] w_sys_tmp8927;
	wire signed [31:0] w_sys_tmp8932;
	wire signed [31:0] w_sys_tmp8933;
	wire signed [31:0] w_sys_tmp8938;
	wire signed [31:0] w_sys_tmp8939;
	wire signed [31:0] w_sys_tmp8944;
	wire signed [31:0] w_sys_tmp8945;
	wire signed [31:0] w_sys_tmp8950;
	wire signed [31:0] w_sys_tmp8951;
	wire signed [31:0] w_sys_tmp8956;
	wire signed [31:0] w_sys_tmp8957;
	wire signed [31:0] w_sys_tmp8962;
	wire signed [31:0] w_sys_tmp8963;
	wire signed [31:0] w_sys_tmp8968;
	wire signed [31:0] w_sys_tmp8969;
	wire signed [31:0] w_sys_tmp8974;
	wire signed [31:0] w_sys_tmp8975;
	wire signed [31:0] w_sys_tmp8980;
	wire signed [31:0] w_sys_tmp8981;
	wire signed [31:0] w_sys_tmp8986;
	wire signed [31:0] w_sys_tmp8987;
	wire signed [31:0] w_sys_tmp8992;
	wire signed [31:0] w_sys_tmp8993;
	wire signed [31:0] w_sys_tmp8998;
	wire signed [31:0] w_sys_tmp8999;
	wire signed [31:0] w_sys_tmp9004;
	wire signed [31:0] w_sys_tmp9005;
	wire signed [31:0] w_sys_tmp9010;
	wire signed [31:0] w_sys_tmp9011;
	wire signed [31:0] w_sys_tmp9016;
	wire signed [31:0] w_sys_tmp9017;
	wire signed [31:0] w_sys_tmp9034;
	wire signed [31:0] w_sys_tmp9035;
	wire signed [31:0] w_sys_tmp9040;
	wire signed [31:0] w_sys_tmp9041;
	wire signed [31:0] w_sys_tmp9046;
	wire signed [31:0] w_sys_tmp9047;
	wire signed [31:0] w_sys_tmp9052;
	wire signed [31:0] w_sys_tmp9053;
	wire signed [31:0] w_sys_tmp9058;
	wire signed [31:0] w_sys_tmp9059;
	wire signed [31:0] w_sys_tmp9064;
	wire signed [31:0] w_sys_tmp9065;
	wire signed [31:0] w_sys_tmp9070;
	wire signed [31:0] w_sys_tmp9071;
	wire signed [31:0] w_sys_tmp9076;
	wire signed [31:0] w_sys_tmp9077;
	wire signed [31:0] w_sys_tmp9082;
	wire signed [31:0] w_sys_tmp9083;
	wire signed [31:0] w_sys_tmp9088;
	wire signed [31:0] w_sys_tmp9089;
	wire signed [31:0] w_sys_tmp9094;
	wire signed [31:0] w_sys_tmp9095;
	wire signed [31:0] w_sys_tmp9100;
	wire signed [31:0] w_sys_tmp9101;
	wire signed [31:0] w_sys_tmp9106;
	wire signed [31:0] w_sys_tmp9107;
	wire signed [31:0] w_sys_tmp9112;
	wire signed [31:0] w_sys_tmp9113;
	wire signed [31:0] w_sys_tmp9118;
	wire signed [31:0] w_sys_tmp9119;
	wire signed [31:0] w_sys_tmp9124;
	wire signed [31:0] w_sys_tmp9125;
	wire signed [31:0] w_sys_tmp9130;
	wire signed [31:0] w_sys_tmp9131;
	wire signed [31:0] w_sys_tmp9136;
	wire signed [31:0] w_sys_tmp9137;
	wire signed [31:0] w_sys_tmp9142;
	wire signed [31:0] w_sys_tmp9143;
	wire signed [31:0] w_sys_tmp9148;
	wire signed [31:0] w_sys_tmp9149;
	wire signed [31:0] w_sys_tmp9166;
	wire signed [31:0] w_sys_tmp9167;
	wire signed [31:0] w_sys_tmp9172;
	wire signed [31:0] w_sys_tmp9173;
	wire signed [31:0] w_sys_tmp9178;
	wire signed [31:0] w_sys_tmp9179;
	wire signed [31:0] w_sys_tmp9184;
	wire signed [31:0] w_sys_tmp9185;
	wire signed [31:0] w_sys_tmp9190;
	wire signed [31:0] w_sys_tmp9191;
	wire signed [31:0] w_sys_tmp9196;
	wire signed [31:0] w_sys_tmp9197;
	wire signed [31:0] w_sys_tmp9202;
	wire signed [31:0] w_sys_tmp9203;
	wire signed [31:0] w_sys_tmp9208;
	wire signed [31:0] w_sys_tmp9209;
	wire signed [31:0] w_sys_tmp9214;
	wire signed [31:0] w_sys_tmp9215;
	wire signed [31:0] w_sys_tmp9220;
	wire signed [31:0] w_sys_tmp9221;
	wire signed [31:0] w_sys_tmp9226;
	wire signed [31:0] w_sys_tmp9227;
	wire signed [31:0] w_sys_tmp9232;
	wire signed [31:0] w_sys_tmp9233;
	wire signed [31:0] w_sys_tmp9238;
	wire signed [31:0] w_sys_tmp9239;
	wire signed [31:0] w_sys_tmp9244;
	wire signed [31:0] w_sys_tmp9245;
	wire signed [31:0] w_sys_tmp9250;
	wire signed [31:0] w_sys_tmp9251;
	wire signed [31:0] w_sys_tmp9256;
	wire signed [31:0] w_sys_tmp9257;
	wire signed [31:0] w_sys_tmp9262;
	wire signed [31:0] w_sys_tmp9263;
	wire signed [31:0] w_sys_tmp9268;
	wire signed [31:0] w_sys_tmp9269;
	wire signed [31:0] w_sys_tmp9274;
	wire signed [31:0] w_sys_tmp9275;
	wire signed [31:0] w_sys_tmp9280;
	wire signed [31:0] w_sys_tmp9281;
	wire signed [31:0] w_sys_tmp9298;
	wire signed [31:0] w_sys_tmp9299;
	wire signed [31:0] w_sys_tmp9304;
	wire signed [31:0] w_sys_tmp9305;
	wire signed [31:0] w_sys_tmp9310;
	wire signed [31:0] w_sys_tmp9311;
	wire signed [31:0] w_sys_tmp9316;
	wire signed [31:0] w_sys_tmp9317;
	wire signed [31:0] w_sys_tmp9322;
	wire signed [31:0] w_sys_tmp9323;
	wire signed [31:0] w_sys_tmp9328;
	wire signed [31:0] w_sys_tmp9329;
	wire signed [31:0] w_sys_tmp9334;
	wire signed [31:0] w_sys_tmp9335;
	wire signed [31:0] w_sys_tmp9340;
	wire signed [31:0] w_sys_tmp9341;
	wire signed [31:0] w_sys_tmp9346;
	wire signed [31:0] w_sys_tmp9347;
	wire signed [31:0] w_sys_tmp9352;
	wire signed [31:0] w_sys_tmp9353;
	wire signed [31:0] w_sys_tmp9358;
	wire signed [31:0] w_sys_tmp9359;
	wire signed [31:0] w_sys_tmp9364;
	wire signed [31:0] w_sys_tmp9365;
	wire signed [31:0] w_sys_tmp9370;
	wire signed [31:0] w_sys_tmp9371;
	wire signed [31:0] w_sys_tmp9376;
	wire signed [31:0] w_sys_tmp9377;
	wire signed [31:0] w_sys_tmp9382;
	wire signed [31:0] w_sys_tmp9383;
	wire signed [31:0] w_sys_tmp9388;
	wire signed [31:0] w_sys_tmp9389;
	wire signed [31:0] w_sys_tmp9394;
	wire signed [31:0] w_sys_tmp9395;
	wire signed [31:0] w_sys_tmp9400;
	wire signed [31:0] w_sys_tmp9401;
	wire signed [31:0] w_sys_tmp9406;
	wire signed [31:0] w_sys_tmp9407;
	wire signed [31:0] w_sys_tmp9412;
	wire signed [31:0] w_sys_tmp9413;
	wire signed [31:0] w_sys_tmp9418;
	wire signed [31:0] w_sys_tmp9419;
	wire signed [31:0] w_sys_tmp9424;
	wire signed [31:0] w_sys_tmp9425;
	wire signed [31:0] w_sys_tmp9430;
	wire signed [31:0] w_sys_tmp9431;
	wire signed [31:0] w_sys_tmp9436;
	wire signed [31:0] w_sys_tmp9437;
	wire signed [31:0] w_sys_tmp9442;
	wire signed [31:0] w_sys_tmp9443;
	wire signed [31:0] w_sys_tmp9448;
	wire signed [31:0] w_sys_tmp9449;
	wire signed [31:0] w_sys_tmp9454;
	wire signed [31:0] w_sys_tmp9455;
	wire signed [31:0] w_sys_tmp9460;
	wire signed [31:0] w_sys_tmp9461;
	wire signed [31:0] w_sys_tmp9466;
	wire signed [31:0] w_sys_tmp9467;
	wire signed [31:0] w_sys_tmp9472;
	wire signed [31:0] w_sys_tmp9473;
	wire signed [31:0] w_sys_tmp9478;
	wire signed [31:0] w_sys_tmp9479;
	wire signed [31:0] w_sys_tmp9484;
	wire signed [31:0] w_sys_tmp9485;
	wire signed [31:0] w_sys_tmp9490;
	wire signed [31:0] w_sys_tmp9491;
	wire signed [31:0] w_sys_tmp9496;
	wire signed [31:0] w_sys_tmp9497;
	wire signed [31:0] w_sys_tmp9502;
	wire signed [31:0] w_sys_tmp9503;
	wire signed [31:0] w_sys_tmp9508;
	wire signed [31:0] w_sys_tmp9509;
	wire signed [31:0] w_sys_tmp9514;
	wire signed [31:0] w_sys_tmp9515;
	wire signed [31:0] w_sys_tmp9520;
	wire signed [31:0] w_sys_tmp9521;
	wire signed [31:0] w_sys_tmp9526;
	wire signed [31:0] w_sys_tmp9527;
	wire signed [31:0] w_sys_tmp9532;
	wire signed [31:0] w_sys_tmp9533;
	wire signed [31:0] w_sys_tmp9538;
	wire signed [31:0] w_sys_tmp9539;
	wire signed [31:0] w_sys_tmp9556;
	wire signed [31:0] w_sys_tmp9557;
	wire signed [31:0] w_sys_tmp9562;
	wire signed [31:0] w_sys_tmp9563;
	wire signed [31:0] w_sys_tmp9568;
	wire signed [31:0] w_sys_tmp9569;
	wire signed [31:0] w_sys_tmp9574;
	wire signed [31:0] w_sys_tmp9575;
	wire signed [31:0] w_sys_tmp9580;
	wire signed [31:0] w_sys_tmp9581;
	wire signed [31:0] w_sys_tmp9586;
	wire signed [31:0] w_sys_tmp9587;
	wire signed [31:0] w_sys_tmp9592;
	wire signed [31:0] w_sys_tmp9593;
	wire signed [31:0] w_sys_tmp9598;
	wire signed [31:0] w_sys_tmp9599;
	wire signed [31:0] w_sys_tmp9604;
	wire signed [31:0] w_sys_tmp9605;
	wire signed [31:0] w_sys_tmp9610;
	wire signed [31:0] w_sys_tmp9611;
	wire signed [31:0] w_sys_tmp9616;
	wire signed [31:0] w_sys_tmp9617;
	wire signed [31:0] w_sys_tmp9622;
	wire signed [31:0] w_sys_tmp9623;
	wire signed [31:0] w_sys_tmp9628;
	wire signed [31:0] w_sys_tmp9629;
	wire signed [31:0] w_sys_tmp9634;
	wire signed [31:0] w_sys_tmp9635;
	wire signed [31:0] w_sys_tmp9640;
	wire signed [31:0] w_sys_tmp9641;
	wire signed [31:0] w_sys_tmp9646;
	wire signed [31:0] w_sys_tmp9647;
	wire signed [31:0] w_sys_tmp9652;
	wire signed [31:0] w_sys_tmp9653;
	wire signed [31:0] w_sys_tmp9658;
	wire signed [31:0] w_sys_tmp9659;
	wire signed [31:0] w_sys_tmp9664;
	wire signed [31:0] w_sys_tmp9665;
	wire signed [31:0] w_sys_tmp9670;
	wire signed [31:0] w_sys_tmp9671;
	wire signed [31:0] w_sys_tmp9688;
	wire signed [31:0] w_sys_tmp9689;
	wire signed [31:0] w_sys_tmp9694;
	wire signed [31:0] w_sys_tmp9695;
	wire signed [31:0] w_sys_tmp9700;
	wire signed [31:0] w_sys_tmp9701;
	wire signed [31:0] w_sys_tmp9706;
	wire signed [31:0] w_sys_tmp9707;
	wire signed [31:0] w_sys_tmp9712;
	wire signed [31:0] w_sys_tmp9713;
	wire signed [31:0] w_sys_tmp9718;
	wire signed [31:0] w_sys_tmp9719;
	wire signed [31:0] w_sys_tmp9724;
	wire signed [31:0] w_sys_tmp9725;
	wire signed [31:0] w_sys_tmp9730;
	wire signed [31:0] w_sys_tmp9731;
	wire signed [31:0] w_sys_tmp9736;
	wire signed [31:0] w_sys_tmp9737;
	wire signed [31:0] w_sys_tmp9742;
	wire signed [31:0] w_sys_tmp9743;
	wire signed [31:0] w_sys_tmp9748;
	wire signed [31:0] w_sys_tmp9749;
	wire signed [31:0] w_sys_tmp9754;
	wire signed [31:0] w_sys_tmp9755;
	wire signed [31:0] w_sys_tmp9760;
	wire signed [31:0] w_sys_tmp9761;
	wire signed [31:0] w_sys_tmp9766;
	wire signed [31:0] w_sys_tmp9767;
	wire signed [31:0] w_sys_tmp9772;
	wire signed [31:0] w_sys_tmp9773;
	wire signed [31:0] w_sys_tmp9778;
	wire signed [31:0] w_sys_tmp9779;
	wire signed [31:0] w_sys_tmp9784;
	wire signed [31:0] w_sys_tmp9785;
	wire signed [31:0] w_sys_tmp9790;
	wire signed [31:0] w_sys_tmp9791;
	wire signed [31:0] w_sys_tmp9796;
	wire signed [31:0] w_sys_tmp9797;
	wire signed [31:0] w_sys_tmp9802;
	wire signed [31:0] w_sys_tmp9803;
	wire signed [31:0] w_sys_tmp9820;
	wire signed [31:0] w_sys_tmp9821;
	wire signed [31:0] w_sys_tmp9826;
	wire signed [31:0] w_sys_tmp9827;
	wire signed [31:0] w_sys_tmp9832;
	wire signed [31:0] w_sys_tmp9833;
	wire signed [31:0] w_sys_tmp9838;
	wire signed [31:0] w_sys_tmp9839;
	wire signed [31:0] w_sys_tmp9844;
	wire signed [31:0] w_sys_tmp9845;
	wire signed [31:0] w_sys_tmp9850;
	wire signed [31:0] w_sys_tmp9851;
	wire signed [31:0] w_sys_tmp9856;
	wire signed [31:0] w_sys_tmp9857;
	wire signed [31:0] w_sys_tmp9862;
	wire signed [31:0] w_sys_tmp9863;
	wire signed [31:0] w_sys_tmp9868;
	wire signed [31:0] w_sys_tmp9869;
	wire signed [31:0] w_sys_tmp9874;
	wire signed [31:0] w_sys_tmp9875;
	wire signed [31:0] w_sys_tmp9880;
	wire signed [31:0] w_sys_tmp9881;
	wire signed [31:0] w_sys_tmp9886;
	wire signed [31:0] w_sys_tmp9887;
	wire signed [31:0] w_sys_tmp9892;
	wire signed [31:0] w_sys_tmp9893;
	wire signed [31:0] w_sys_tmp9898;
	wire signed [31:0] w_sys_tmp9899;
	wire signed [31:0] w_sys_tmp9904;
	wire signed [31:0] w_sys_tmp9905;
	wire signed [31:0] w_sys_tmp9910;
	wire signed [31:0] w_sys_tmp9911;
	wire signed [31:0] w_sys_tmp9916;
	wire signed [31:0] w_sys_tmp9917;
	wire signed [31:0] w_sys_tmp9922;
	wire signed [31:0] w_sys_tmp9923;
	wire signed [31:0] w_sys_tmp9928;
	wire signed [31:0] w_sys_tmp9929;
	wire signed [31:0] w_sys_tmp9934;
	wire signed [31:0] w_sys_tmp9935;
	wire signed [31:0] w_sys_tmp9952;
	wire signed [31:0] w_sys_tmp9953;
	wire signed [31:0] w_sys_tmp9958;
	wire signed [31:0] w_sys_tmp9959;
	wire signed [31:0] w_sys_tmp9964;
	wire signed [31:0] w_sys_tmp9965;
	wire signed [31:0] w_sys_tmp9970;
	wire signed [31:0] w_sys_tmp9971;
	wire signed [31:0] w_sys_tmp9976;
	wire signed [31:0] w_sys_tmp9977;
	wire signed [31:0] w_sys_tmp9982;
	wire signed [31:0] w_sys_tmp9983;
	wire signed [31:0] w_sys_tmp9988;
	wire signed [31:0] w_sys_tmp9989;
	wire signed [31:0] w_sys_tmp9994;
	wire signed [31:0] w_sys_tmp9995;
	wire signed [31:0] w_sys_tmp10000;
	wire signed [31:0] w_sys_tmp10001;
	wire signed [31:0] w_sys_tmp10006;
	wire signed [31:0] w_sys_tmp10007;
	wire signed [31:0] w_sys_tmp10012;
	wire signed [31:0] w_sys_tmp10013;
	wire signed [31:0] w_sys_tmp10018;
	wire signed [31:0] w_sys_tmp10019;
	wire signed [31:0] w_sys_tmp10024;
	wire signed [31:0] w_sys_tmp10025;
	wire signed [31:0] w_sys_tmp10030;
	wire signed [31:0] w_sys_tmp10031;
	wire signed [31:0] w_sys_tmp10036;
	wire signed [31:0] w_sys_tmp10037;
	wire signed [31:0] w_sys_tmp10042;
	wire signed [31:0] w_sys_tmp10043;
	wire signed [31:0] w_sys_tmp10048;
	wire signed [31:0] w_sys_tmp10049;
	wire signed [31:0] w_sys_tmp10054;
	wire signed [31:0] w_sys_tmp10055;
	wire signed [31:0] w_sys_tmp10060;
	wire signed [31:0] w_sys_tmp10061;
	wire signed [31:0] w_sys_tmp10065;
	wire signed [31:0] w_sys_tmp10066;
	wire               w_sys_tmp10067;
	wire               w_sys_tmp10068;
	wire signed [31:0] w_sys_tmp10069;
	wire signed [31:0] w_sys_tmp10072;
	wire signed [31:0] w_sys_tmp10073;
	wire        [31:0] w_sys_tmp10074;
	wire signed [31:0] w_sys_tmp10078;
	wire signed [31:0] w_sys_tmp10079;
	wire signed [31:0] w_sys_tmp10084;
	wire signed [31:0] w_sys_tmp10085;
	wire signed [31:0] w_sys_tmp10090;
	wire signed [31:0] w_sys_tmp10091;
	wire signed [31:0] w_sys_tmp10096;
	wire signed [31:0] w_sys_tmp10097;
	wire signed [31:0] w_sys_tmp10102;
	wire signed [31:0] w_sys_tmp10103;
	wire signed [31:0] w_sys_tmp10108;
	wire signed [31:0] w_sys_tmp10109;
	wire signed [31:0] w_sys_tmp10114;
	wire signed [31:0] w_sys_tmp10115;
	wire signed [31:0] w_sys_tmp10120;
	wire signed [31:0] w_sys_tmp10121;
	wire signed [31:0] w_sys_tmp10126;
	wire signed [31:0] w_sys_tmp10127;
	wire signed [31:0] w_sys_tmp10132;
	wire signed [31:0] w_sys_tmp10133;
	wire signed [31:0] w_sys_tmp10138;
	wire signed [31:0] w_sys_tmp10139;
	wire signed [31:0] w_sys_tmp10144;
	wire signed [31:0] w_sys_tmp10145;
	wire signed [31:0] w_sys_tmp10150;
	wire signed [31:0] w_sys_tmp10151;
	wire signed [31:0] w_sys_tmp10156;
	wire signed [31:0] w_sys_tmp10157;
	wire signed [31:0] w_sys_tmp10162;
	wire signed [31:0] w_sys_tmp10163;
	wire signed [31:0] w_sys_tmp10168;
	wire signed [31:0] w_sys_tmp10169;
	wire signed [31:0] w_sys_tmp10174;
	wire signed [31:0] w_sys_tmp10175;
	wire signed [31:0] w_sys_tmp10180;
	wire signed [31:0] w_sys_tmp10181;
	wire signed [31:0] w_sys_tmp10186;
	wire signed [31:0] w_sys_tmp10187;
	wire signed [31:0] w_sys_tmp10192;
	wire signed [31:0] w_sys_tmp10193;
	wire signed [31:0] w_sys_tmp10198;
	wire signed [31:0] w_sys_tmp10199;
	wire signed [31:0] w_sys_tmp10216;
	wire signed [31:0] w_sys_tmp10217;
	wire signed [31:0] w_sys_tmp10222;
	wire signed [31:0] w_sys_tmp10223;
	wire signed [31:0] w_sys_tmp10228;
	wire signed [31:0] w_sys_tmp10229;
	wire signed [31:0] w_sys_tmp10234;
	wire signed [31:0] w_sys_tmp10235;
	wire signed [31:0] w_sys_tmp10240;
	wire signed [31:0] w_sys_tmp10241;
	wire signed [31:0] w_sys_tmp10246;
	wire signed [31:0] w_sys_tmp10247;
	wire signed [31:0] w_sys_tmp10252;
	wire signed [31:0] w_sys_tmp10253;
	wire signed [31:0] w_sys_tmp10258;
	wire signed [31:0] w_sys_tmp10259;
	wire signed [31:0] w_sys_tmp10264;
	wire signed [31:0] w_sys_tmp10265;
	wire signed [31:0] w_sys_tmp10270;
	wire signed [31:0] w_sys_tmp10271;
	wire signed [31:0] w_sys_tmp10276;
	wire signed [31:0] w_sys_tmp10277;
	wire signed [31:0] w_sys_tmp10282;
	wire signed [31:0] w_sys_tmp10283;
	wire signed [31:0] w_sys_tmp10288;
	wire signed [31:0] w_sys_tmp10289;
	wire signed [31:0] w_sys_tmp10294;
	wire signed [31:0] w_sys_tmp10295;
	wire signed [31:0] w_sys_tmp10300;
	wire signed [31:0] w_sys_tmp10301;
	wire signed [31:0] w_sys_tmp10306;
	wire signed [31:0] w_sys_tmp10307;
	wire signed [31:0] w_sys_tmp10312;
	wire signed [31:0] w_sys_tmp10313;
	wire signed [31:0] w_sys_tmp10318;
	wire signed [31:0] w_sys_tmp10319;
	wire signed [31:0] w_sys_tmp10324;
	wire signed [31:0] w_sys_tmp10325;
	wire signed [31:0] w_sys_tmp10330;
	wire signed [31:0] w_sys_tmp10331;
	wire signed [31:0] w_sys_tmp10348;
	wire signed [31:0] w_sys_tmp10349;
	wire signed [31:0] w_sys_tmp10354;
	wire signed [31:0] w_sys_tmp10355;
	wire signed [31:0] w_sys_tmp10360;
	wire signed [31:0] w_sys_tmp10361;
	wire signed [31:0] w_sys_tmp10366;
	wire signed [31:0] w_sys_tmp10367;
	wire signed [31:0] w_sys_tmp10372;
	wire signed [31:0] w_sys_tmp10373;
	wire signed [31:0] w_sys_tmp10378;
	wire signed [31:0] w_sys_tmp10379;
	wire signed [31:0] w_sys_tmp10384;
	wire signed [31:0] w_sys_tmp10385;
	wire signed [31:0] w_sys_tmp10390;
	wire signed [31:0] w_sys_tmp10391;
	wire signed [31:0] w_sys_tmp10396;
	wire signed [31:0] w_sys_tmp10397;
	wire signed [31:0] w_sys_tmp10402;
	wire signed [31:0] w_sys_tmp10403;
	wire signed [31:0] w_sys_tmp10408;
	wire signed [31:0] w_sys_tmp10409;
	wire signed [31:0] w_sys_tmp10414;
	wire signed [31:0] w_sys_tmp10415;
	wire signed [31:0] w_sys_tmp10420;
	wire signed [31:0] w_sys_tmp10421;
	wire signed [31:0] w_sys_tmp10426;
	wire signed [31:0] w_sys_tmp10427;
	wire signed [31:0] w_sys_tmp10432;
	wire signed [31:0] w_sys_tmp10433;
	wire signed [31:0] w_sys_tmp10438;
	wire signed [31:0] w_sys_tmp10439;
	wire signed [31:0] w_sys_tmp10444;
	wire signed [31:0] w_sys_tmp10445;
	wire signed [31:0] w_sys_tmp10450;
	wire signed [31:0] w_sys_tmp10451;
	wire signed [31:0] w_sys_tmp10456;
	wire signed [31:0] w_sys_tmp10457;
	wire signed [31:0] w_sys_tmp10462;
	wire signed [31:0] w_sys_tmp10463;
	wire signed [31:0] w_sys_tmp10480;
	wire signed [31:0] w_sys_tmp10481;
	wire signed [31:0] w_sys_tmp10486;
	wire signed [31:0] w_sys_tmp10487;
	wire signed [31:0] w_sys_tmp10492;
	wire signed [31:0] w_sys_tmp10493;
	wire signed [31:0] w_sys_tmp10498;
	wire signed [31:0] w_sys_tmp10499;
	wire signed [31:0] w_sys_tmp10504;
	wire signed [31:0] w_sys_tmp10505;
	wire signed [31:0] w_sys_tmp10510;
	wire signed [31:0] w_sys_tmp10511;
	wire signed [31:0] w_sys_tmp10516;
	wire signed [31:0] w_sys_tmp10517;
	wire signed [31:0] w_sys_tmp10522;
	wire signed [31:0] w_sys_tmp10523;
	wire signed [31:0] w_sys_tmp10528;
	wire signed [31:0] w_sys_tmp10529;
	wire signed [31:0] w_sys_tmp10534;
	wire signed [31:0] w_sys_tmp10535;
	wire signed [31:0] w_sys_tmp10540;
	wire signed [31:0] w_sys_tmp10541;
	wire signed [31:0] w_sys_tmp10546;
	wire signed [31:0] w_sys_tmp10547;
	wire signed [31:0] w_sys_tmp10552;
	wire signed [31:0] w_sys_tmp10553;
	wire signed [31:0] w_sys_tmp10558;
	wire signed [31:0] w_sys_tmp10559;
	wire signed [31:0] w_sys_tmp10564;
	wire signed [31:0] w_sys_tmp10565;
	wire signed [31:0] w_sys_tmp10570;
	wire signed [31:0] w_sys_tmp10571;
	wire signed [31:0] w_sys_tmp10576;
	wire signed [31:0] w_sys_tmp10577;
	wire signed [31:0] w_sys_tmp10582;
	wire signed [31:0] w_sys_tmp10583;
	wire signed [31:0] w_sys_tmp10588;
	wire signed [31:0] w_sys_tmp10589;
	wire signed [31:0] w_sys_tmp10594;
	wire signed [31:0] w_sys_tmp10595;
	wire signed [31:0] w_sys_tmp10612;
	wire signed [31:0] w_sys_tmp10613;
	wire signed [31:0] w_sys_tmp10618;
	wire signed [31:0] w_sys_tmp10619;
	wire signed [31:0] w_sys_tmp10624;
	wire signed [31:0] w_sys_tmp10625;
	wire signed [31:0] w_sys_tmp10630;
	wire signed [31:0] w_sys_tmp10631;
	wire signed [31:0] w_sys_tmp10636;
	wire signed [31:0] w_sys_tmp10637;
	wire signed [31:0] w_sys_tmp10642;
	wire signed [31:0] w_sys_tmp10643;
	wire signed [31:0] w_sys_tmp10648;
	wire signed [31:0] w_sys_tmp10649;
	wire signed [31:0] w_sys_tmp10654;
	wire signed [31:0] w_sys_tmp10655;
	wire signed [31:0] w_sys_tmp10660;
	wire signed [31:0] w_sys_tmp10661;
	wire signed [31:0] w_sys_tmp10666;
	wire signed [31:0] w_sys_tmp10667;
	wire signed [31:0] w_sys_tmp10672;
	wire signed [31:0] w_sys_tmp10673;
	wire signed [31:0] w_sys_tmp10678;
	wire signed [31:0] w_sys_tmp10679;
	wire signed [31:0] w_sys_tmp10684;
	wire signed [31:0] w_sys_tmp10685;
	wire signed [31:0] w_sys_tmp10690;
	wire signed [31:0] w_sys_tmp10691;
	wire signed [31:0] w_sys_tmp10696;
	wire signed [31:0] w_sys_tmp10697;
	wire signed [31:0] w_sys_tmp10702;
	wire signed [31:0] w_sys_tmp10703;
	wire signed [31:0] w_sys_tmp10708;
	wire signed [31:0] w_sys_tmp10709;
	wire signed [31:0] w_sys_tmp10714;
	wire signed [31:0] w_sys_tmp10715;
	wire signed [31:0] w_sys_tmp10720;
	wire signed [31:0] w_sys_tmp10721;
	wire signed [31:0] w_sys_tmp10725;
	wire signed [31:0] w_sys_tmp10726;
	wire               w_sys_tmp10727;
	wire               w_sys_tmp10728;
	wire signed [31:0] w_sys_tmp10729;
	wire signed [31:0] w_sys_tmp10732;
	wire signed [31:0] w_sys_tmp10733;
	wire        [31:0] w_sys_tmp10734;
	wire signed [31:0] w_sys_tmp10738;
	wire signed [31:0] w_sys_tmp10739;
	wire signed [31:0] w_sys_tmp10744;
	wire signed [31:0] w_sys_tmp10745;
	wire signed [31:0] w_sys_tmp10750;
	wire signed [31:0] w_sys_tmp10751;
	wire signed [31:0] w_sys_tmp10756;
	wire signed [31:0] w_sys_tmp10757;
	wire signed [31:0] w_sys_tmp10762;
	wire signed [31:0] w_sys_tmp10763;
	wire signed [31:0] w_sys_tmp10768;
	wire signed [31:0] w_sys_tmp10769;
	wire signed [31:0] w_sys_tmp10774;
	wire signed [31:0] w_sys_tmp10775;
	wire signed [31:0] w_sys_tmp10780;
	wire signed [31:0] w_sys_tmp10781;
	wire signed [31:0] w_sys_tmp10786;
	wire signed [31:0] w_sys_tmp10787;
	wire signed [31:0] w_sys_tmp10792;
	wire signed [31:0] w_sys_tmp10793;
	wire signed [31:0] w_sys_tmp10798;
	wire signed [31:0] w_sys_tmp10799;
	wire signed [31:0] w_sys_tmp10804;
	wire signed [31:0] w_sys_tmp10805;
	wire signed [31:0] w_sys_tmp10810;
	wire signed [31:0] w_sys_tmp10811;
	wire signed [31:0] w_sys_tmp10816;
	wire signed [31:0] w_sys_tmp10817;
	wire signed [31:0] w_sys_tmp10822;
	wire signed [31:0] w_sys_tmp10823;
	wire signed [31:0] w_sys_tmp10828;
	wire signed [31:0] w_sys_tmp10829;
	wire signed [31:0] w_sys_tmp10834;
	wire signed [31:0] w_sys_tmp10835;
	wire signed [31:0] w_sys_tmp10840;
	wire signed [31:0] w_sys_tmp10841;
	wire signed [31:0] w_sys_tmp10846;
	wire signed [31:0] w_sys_tmp10847;
	wire signed [31:0] w_sys_tmp10922;
	wire signed [31:0] w_sys_tmp10923;
	wire signed [31:0] w_sys_tmp10927;
	wire signed [31:0] w_sys_tmp10928;
	wire signed [31:0] w_sys_tmp10932;
	wire signed [31:0] w_sys_tmp10933;
	wire signed [31:0] w_sys_tmp10937;
	wire signed [31:0] w_sys_tmp10938;
	wire signed [31:0] w_sys_tmp10942;
	wire signed [31:0] w_sys_tmp10943;
	wire signed [31:0] w_sys_tmp10947;
	wire signed [31:0] w_sys_tmp10948;
	wire signed [31:0] w_sys_tmp10952;
	wire signed [31:0] w_sys_tmp10953;
	wire signed [31:0] w_sys_tmp10957;
	wire signed [31:0] w_sys_tmp10958;
	wire signed [31:0] w_sys_tmp10962;
	wire signed [31:0] w_sys_tmp10963;
	wire signed [31:0] w_sys_tmp10967;
	wire signed [31:0] w_sys_tmp10968;
	wire signed [31:0] w_sys_tmp10972;
	wire signed [31:0] w_sys_tmp10973;
	wire signed [31:0] w_sys_tmp10977;
	wire signed [31:0] w_sys_tmp10978;
	wire signed [31:0] w_sys_tmp10982;
	wire signed [31:0] w_sys_tmp10983;
	wire signed [31:0] w_sys_tmp10987;
	wire signed [31:0] w_sys_tmp10988;
	wire signed [31:0] w_sys_tmp10992;
	wire signed [31:0] w_sys_tmp10993;
	wire signed [31:0] w_sys_tmp10997;
	wire signed [31:0] w_sys_tmp10998;
	wire signed [31:0] w_sys_tmp11002;
	wire signed [31:0] w_sys_tmp11003;
	wire signed [31:0] w_sys_tmp11007;
	wire signed [31:0] w_sys_tmp11008;
	wire signed [31:0] w_sys_tmp11012;
	wire signed [31:0] w_sys_tmp11013;
	wire signed [31:0] w_sys_tmp11017;
	wire signed [31:0] w_sys_tmp11018;
	wire signed [31:0] w_sys_tmp11162;
	wire signed [31:0] w_sys_tmp11163;
	wire signed [31:0] w_sys_tmp11167;
	wire signed [31:0] w_sys_tmp11168;
	wire signed [31:0] w_sys_tmp11172;
	wire signed [31:0] w_sys_tmp11173;
	wire signed [31:0] w_sys_tmp11177;
	wire signed [31:0] w_sys_tmp11178;
	wire signed [31:0] w_sys_tmp11182;
	wire signed [31:0] w_sys_tmp11183;
	wire signed [31:0] w_sys_tmp11187;
	wire signed [31:0] w_sys_tmp11188;
	wire signed [31:0] w_sys_tmp11192;
	wire signed [31:0] w_sys_tmp11193;
	wire signed [31:0] w_sys_tmp11197;
	wire signed [31:0] w_sys_tmp11198;
	wire signed [31:0] w_sys_tmp11202;
	wire signed [31:0] w_sys_tmp11203;
	wire signed [31:0] w_sys_tmp11207;
	wire signed [31:0] w_sys_tmp11208;
	wire signed [31:0] w_sys_tmp11212;
	wire signed [31:0] w_sys_tmp11213;
	wire signed [31:0] w_sys_tmp11217;
	wire signed [31:0] w_sys_tmp11218;
	wire signed [31:0] w_sys_tmp11222;
	wire signed [31:0] w_sys_tmp11223;
	wire signed [31:0] w_sys_tmp11227;
	wire signed [31:0] w_sys_tmp11228;
	wire signed [31:0] w_sys_tmp11232;
	wire signed [31:0] w_sys_tmp11233;
	wire signed [31:0] w_sys_tmp11237;
	wire signed [31:0] w_sys_tmp11238;
	wire signed [31:0] w_sys_tmp11242;
	wire signed [31:0] w_sys_tmp11243;
	wire signed [31:0] w_sys_tmp11247;
	wire signed [31:0] w_sys_tmp11248;
	wire signed [31:0] w_sys_tmp11252;
	wire signed [31:0] w_sys_tmp11253;
	wire signed [31:0] w_sys_tmp11257;
	wire signed [31:0] w_sys_tmp11258;
	wire signed [31:0] w_sys_tmp11267;
	wire signed [31:0] w_sys_tmp11268;
	wire signed [31:0] w_sys_tmp11272;
	wire signed [31:0] w_sys_tmp11273;
	wire signed [31:0] w_sys_tmp11277;
	wire signed [31:0] w_sys_tmp11278;
	wire signed [31:0] w_sys_tmp11282;
	wire signed [31:0] w_sys_tmp11283;
	wire signed [31:0] w_sys_tmp11287;
	wire signed [31:0] w_sys_tmp11288;
	wire signed [31:0] w_sys_tmp11292;
	wire signed [31:0] w_sys_tmp11293;
	wire signed [31:0] w_sys_tmp11297;
	wire signed [31:0] w_sys_tmp11298;
	wire signed [31:0] w_sys_tmp11302;
	wire signed [31:0] w_sys_tmp11303;
	wire signed [31:0] w_sys_tmp11307;
	wire signed [31:0] w_sys_tmp11308;
	wire signed [31:0] w_sys_tmp11312;
	wire signed [31:0] w_sys_tmp11313;
	wire signed [31:0] w_sys_tmp11317;
	wire signed [31:0] w_sys_tmp11318;
	wire signed [31:0] w_sys_tmp11322;
	wire signed [31:0] w_sys_tmp11323;
	wire signed [31:0] w_sys_tmp11327;
	wire signed [31:0] w_sys_tmp11328;
	wire signed [31:0] w_sys_tmp11332;
	wire signed [31:0] w_sys_tmp11333;
	wire signed [31:0] w_sys_tmp11337;
	wire signed [31:0] w_sys_tmp11338;
	wire signed [31:0] w_sys_tmp11342;
	wire signed [31:0] w_sys_tmp11343;
	wire signed [31:0] w_sys_tmp11347;
	wire signed [31:0] w_sys_tmp11348;
	wire signed [31:0] w_sys_tmp11352;
	wire signed [31:0] w_sys_tmp11353;
	wire signed [31:0] w_sys_tmp11357;
	wire signed [31:0] w_sys_tmp11358;
	wire signed [31:0] w_sys_tmp11362;
	wire signed [31:0] w_sys_tmp11363;
	wire signed [31:0] w_sys_tmp11372;
	wire signed [31:0] w_sys_tmp11373;
	wire signed [31:0] w_sys_tmp11377;
	wire signed [31:0] w_sys_tmp11378;
	wire signed [31:0] w_sys_tmp11382;
	wire signed [31:0] w_sys_tmp11383;
	wire signed [31:0] w_sys_tmp11387;
	wire signed [31:0] w_sys_tmp11388;
	wire signed [31:0] w_sys_tmp11392;
	wire signed [31:0] w_sys_tmp11393;
	wire signed [31:0] w_sys_tmp11397;
	wire signed [31:0] w_sys_tmp11398;
	wire signed [31:0] w_sys_tmp11402;
	wire signed [31:0] w_sys_tmp11403;
	wire signed [31:0] w_sys_tmp11407;
	wire signed [31:0] w_sys_tmp11408;
	wire signed [31:0] w_sys_tmp11412;
	wire signed [31:0] w_sys_tmp11413;
	wire signed [31:0] w_sys_tmp11417;
	wire signed [31:0] w_sys_tmp11418;
	wire signed [31:0] w_sys_tmp11422;
	wire signed [31:0] w_sys_tmp11423;
	wire signed [31:0] w_sys_tmp11427;
	wire signed [31:0] w_sys_tmp11428;
	wire signed [31:0] w_sys_tmp11432;
	wire signed [31:0] w_sys_tmp11433;
	wire signed [31:0] w_sys_tmp11437;
	wire signed [31:0] w_sys_tmp11438;
	wire signed [31:0] w_sys_tmp11442;
	wire signed [31:0] w_sys_tmp11443;
	wire signed [31:0] w_sys_tmp11447;
	wire signed [31:0] w_sys_tmp11448;
	wire signed [31:0] w_sys_tmp11452;
	wire signed [31:0] w_sys_tmp11453;
	wire signed [31:0] w_sys_tmp11457;
	wire signed [31:0] w_sys_tmp11458;
	wire signed [31:0] w_sys_tmp11462;
	wire signed [31:0] w_sys_tmp11463;
	wire signed [31:0] w_sys_tmp11467;
	wire signed [31:0] w_sys_tmp11468;
	wire signed [31:0] w_sys_tmp11472;
	wire signed [31:0] w_sys_tmp11473;
	wire signed [31:0] w_sys_tmp11477;
	wire signed [31:0] w_sys_tmp11478;
	wire signed [31:0] w_sys_tmp11482;
	wire signed [31:0] w_sys_tmp11483;
	wire signed [31:0] w_sys_tmp11487;
	wire signed [31:0] w_sys_tmp11488;
	wire signed [31:0] w_sys_tmp11492;
	wire signed [31:0] w_sys_tmp11493;
	wire signed [31:0] w_sys_tmp11497;
	wire signed [31:0] w_sys_tmp11498;
	wire signed [31:0] w_sys_tmp11502;
	wire signed [31:0] w_sys_tmp11503;
	wire signed [31:0] w_sys_tmp11507;
	wire signed [31:0] w_sys_tmp11508;
	wire signed [31:0] w_sys_tmp11512;
	wire signed [31:0] w_sys_tmp11513;
	wire signed [31:0] w_sys_tmp11517;
	wire signed [31:0] w_sys_tmp11518;
	wire signed [31:0] w_sys_tmp11522;
	wire signed [31:0] w_sys_tmp11523;
	wire signed [31:0] w_sys_tmp11527;
	wire signed [31:0] w_sys_tmp11528;
	wire signed [31:0] w_sys_tmp11532;
	wire signed [31:0] w_sys_tmp11533;
	wire signed [31:0] w_sys_tmp11537;
	wire signed [31:0] w_sys_tmp11538;
	wire signed [31:0] w_sys_tmp11542;
	wire signed [31:0] w_sys_tmp11543;
	wire signed [31:0] w_sys_tmp11547;
	wire signed [31:0] w_sys_tmp11548;
	wire signed [31:0] w_sys_tmp11552;
	wire signed [31:0] w_sys_tmp11553;
	wire signed [31:0] w_sys_tmp11557;
	wire signed [31:0] w_sys_tmp11558;
	wire signed [31:0] w_sys_tmp11562;
	wire signed [31:0] w_sys_tmp11563;
	wire signed [31:0] w_sys_tmp11567;
	wire signed [31:0] w_sys_tmp11568;
	wire signed [31:0] w_sys_tmp11572;
	wire signed [31:0] w_sys_tmp11573;
	wire signed [31:0] w_sys_tmp11577;
	wire signed [31:0] w_sys_tmp11578;
	wire signed [31:0] w_sys_tmp11582;
	wire signed [31:0] w_sys_tmp11583;
	wire signed [31:0] w_sys_tmp11587;
	wire signed [31:0] w_sys_tmp11588;
	wire signed [31:0] w_sys_tmp11592;
	wire signed [31:0] w_sys_tmp11593;
	wire signed [31:0] w_sys_tmp11597;
	wire signed [31:0] w_sys_tmp11598;
	wire signed [31:0] w_sys_tmp11602;
	wire signed [31:0] w_sys_tmp11603;
	wire signed [31:0] w_sys_tmp11607;
	wire signed [31:0] w_sys_tmp11608;
	wire signed [31:0] w_sys_tmp11612;
	wire signed [31:0] w_sys_tmp11613;
	wire signed [31:0] w_sys_tmp11617;
	wire signed [31:0] w_sys_tmp11618;
	wire signed [31:0] w_sys_tmp11622;
	wire signed [31:0] w_sys_tmp11623;
	wire signed [31:0] w_sys_tmp11627;
	wire signed [31:0] w_sys_tmp11628;
	wire signed [31:0] w_sys_tmp11632;
	wire signed [31:0] w_sys_tmp11633;
	wire signed [31:0] w_sys_tmp11637;
	wire signed [31:0] w_sys_tmp11638;
	wire signed [31:0] w_sys_tmp11642;
	wire signed [31:0] w_sys_tmp11643;
	wire signed [31:0] w_sys_tmp11647;
	wire signed [31:0] w_sys_tmp11648;
	wire signed [31:0] w_sys_tmp11652;
	wire signed [31:0] w_sys_tmp11653;
	wire signed [31:0] w_sys_tmp11657;
	wire signed [31:0] w_sys_tmp11658;
	wire signed [31:0] w_sys_tmp11662;
	wire signed [31:0] w_sys_tmp11663;
	wire signed [31:0] w_sys_tmp11667;
	wire signed [31:0] w_sys_tmp11668;
	wire signed [31:0] w_sys_tmp11672;
	wire signed [31:0] w_sys_tmp11673;
	wire signed [31:0] w_sys_tmp11677;
	wire signed [31:0] w_sys_tmp11678;
	wire signed [31:0] w_sys_tmp11682;
	wire signed [31:0] w_sys_tmp11683;
	wire signed [31:0] w_sys_tmp11687;
	wire signed [31:0] w_sys_tmp11688;
	wire signed [31:0] w_sys_tmp11692;
	wire signed [31:0] w_sys_tmp11693;
	wire signed [31:0] w_sys_tmp11697;
	wire signed [31:0] w_sys_tmp11698;
	wire signed [31:0] w_sys_tmp11702;
	wire signed [31:0] w_sys_tmp11703;
	wire signed [31:0] w_sys_tmp11707;
	wire signed [31:0] w_sys_tmp11708;
	wire signed [31:0] w_sys_tmp11712;
	wire signed [31:0] w_sys_tmp11713;
	wire signed [31:0] w_sys_tmp11717;
	wire signed [31:0] w_sys_tmp11718;
	wire signed [31:0] w_sys_tmp11722;
	wire signed [31:0] w_sys_tmp11723;
	wire signed [31:0] w_sys_tmp11727;
	wire signed [31:0] w_sys_tmp11728;
	wire signed [31:0] w_sys_tmp11732;
	wire signed [31:0] w_sys_tmp11733;
	wire signed [31:0] w_sys_tmp11737;
	wire signed [31:0] w_sys_tmp11738;
	wire signed [31:0] w_sys_tmp11742;
	wire signed [31:0] w_sys_tmp11743;
	wire signed [31:0] w_sys_tmp11747;
	wire signed [31:0] w_sys_tmp11748;
	wire signed [31:0] w_sys_tmp11752;
	wire signed [31:0] w_sys_tmp11753;
	wire signed [31:0] w_sys_tmp11757;
	wire signed [31:0] w_sys_tmp11758;
	wire signed [31:0] w_sys_tmp11762;
	wire signed [31:0] w_sys_tmp11763;
	wire signed [31:0] w_sys_tmp11767;
	wire signed [31:0] w_sys_tmp11768;
	wire signed [31:0] w_sys_tmp11772;
	wire signed [31:0] w_sys_tmp11773;
	wire signed [31:0] w_sys_tmp11777;
	wire signed [31:0] w_sys_tmp11778;
	wire signed [31:0] w_sys_tmp11782;
	wire signed [31:0] w_sys_tmp11783;
	wire signed [31:0] w_sys_tmp11787;
	wire signed [31:0] w_sys_tmp11788;
	wire signed [31:0] w_sys_tmp11792;
	wire signed [31:0] w_sys_tmp11793;
	wire signed [31:0] w_sys_tmp11797;
	wire signed [31:0] w_sys_tmp11798;
	wire signed [31:0] w_sys_tmp11802;
	wire signed [31:0] w_sys_tmp11803;
	wire signed [31:0] w_sys_tmp11807;
	wire signed [31:0] w_sys_tmp11808;
	wire signed [31:0] w_sys_tmp11812;
	wire signed [31:0] w_sys_tmp11813;
	wire signed [31:0] w_sys_tmp11817;
	wire signed [31:0] w_sys_tmp11818;
	wire signed [31:0] w_sys_tmp11822;
	wire signed [31:0] w_sys_tmp11823;
	wire signed [31:0] w_sys_tmp11827;
	wire signed [31:0] w_sys_tmp11828;
	wire signed [31:0] w_sys_tmp11832;
	wire signed [31:0] w_sys_tmp11833;
	wire signed [31:0] w_sys_tmp11837;
	wire signed [31:0] w_sys_tmp11838;
	wire signed [31:0] w_sys_tmp11842;
	wire signed [31:0] w_sys_tmp11843;
	wire signed [31:0] w_sys_tmp11847;
	wire signed [31:0] w_sys_tmp11848;
	wire signed [31:0] w_sys_tmp11852;
	wire signed [31:0] w_sys_tmp11853;
	wire signed [31:0] w_sys_tmp11857;
	wire signed [31:0] w_sys_tmp11858;
	wire signed [31:0] w_sys_tmp11862;
	wire signed [31:0] w_sys_tmp11863;
	wire signed [31:0] w_sys_tmp11867;
	wire signed [31:0] w_sys_tmp11868;
	wire signed [31:0] w_sys_tmp11872;
	wire signed [31:0] w_sys_tmp11873;
	wire signed [31:0] w_sys_tmp11877;
	wire signed [31:0] w_sys_tmp11878;
	wire signed [31:0] w_sys_tmp11882;
	wire signed [31:0] w_sys_tmp11883;
	wire signed [31:0] w_sys_tmp11887;
	wire signed [31:0] w_sys_tmp11888;
	wire signed [31:0] w_sys_tmp11892;
	wire signed [31:0] w_sys_tmp11893;
	wire signed [31:0] w_sys_tmp11897;
	wire signed [31:0] w_sys_tmp11898;
	wire signed [31:0] w_sys_tmp11902;
	wire signed [31:0] w_sys_tmp11903;
	wire signed [31:0] w_sys_tmp11907;
	wire signed [31:0] w_sys_tmp11908;
	wire signed [31:0] w_sys_tmp11912;
	wire signed [31:0] w_sys_tmp11913;
	wire signed [31:0] w_sys_tmp11917;
	wire signed [31:0] w_sys_tmp11918;
	wire signed [31:0] w_sys_tmp11922;
	wire signed [31:0] w_sys_tmp11923;
	wire signed [31:0] w_sys_tmp11927;
	wire signed [31:0] w_sys_tmp11928;
	wire signed [31:0] w_sys_tmp11932;
	wire signed [31:0] w_sys_tmp11933;
	wire signed [31:0] w_sys_tmp11937;
	wire signed [31:0] w_sys_tmp11938;
	wire signed [31:0] w_sys_tmp11942;
	wire signed [31:0] w_sys_tmp11943;
	wire signed [31:0] w_sys_tmp11947;
	wire signed [31:0] w_sys_tmp11948;
	wire signed [31:0] w_sys_tmp11952;
	wire signed [31:0] w_sys_tmp11953;
	wire signed [31:0] w_sys_tmp11957;
	wire signed [31:0] w_sys_tmp11958;
	wire signed [31:0] w_sys_tmp11962;
	wire signed [31:0] w_sys_tmp11963;
	wire signed [31:0] w_sys_tmp11967;
	wire signed [31:0] w_sys_tmp11968;
	wire signed [31:0] w_sys_tmp11972;
	wire signed [31:0] w_sys_tmp11973;
	wire signed [31:0] w_sys_tmp11977;
	wire signed [31:0] w_sys_tmp11978;
	wire signed [31:0] w_sys_tmp11982;
	wire signed [31:0] w_sys_tmp11983;
	wire signed [31:0] w_sys_tmp11987;
	wire signed [31:0] w_sys_tmp11988;
	wire signed [31:0] w_sys_tmp11992;
	wire signed [31:0] w_sys_tmp11993;
	wire signed [31:0] w_sys_tmp11997;
	wire signed [31:0] w_sys_tmp11998;
	wire signed [31:0] w_sys_tmp12002;
	wire signed [31:0] w_sys_tmp12003;
	wire signed [31:0] w_sys_tmp12007;
	wire signed [31:0] w_sys_tmp12008;
	wire signed [31:0] w_sys_tmp12012;
	wire signed [31:0] w_sys_tmp12013;
	wire signed [31:0] w_sys_tmp12017;
	wire signed [31:0] w_sys_tmp12018;
	wire signed [31:0] w_sys_tmp12022;
	wire signed [31:0] w_sys_tmp12023;
	wire signed [31:0] w_sys_tmp12027;
	wire signed [31:0] w_sys_tmp12028;
	wire signed [31:0] w_sys_tmp12032;
	wire signed [31:0] w_sys_tmp12033;
	wire signed [31:0] w_sys_tmp12037;
	wire signed [31:0] w_sys_tmp12038;
	wire signed [31:0] w_sys_tmp12042;
	wire signed [31:0] w_sys_tmp12043;
	wire signed [31:0] w_sys_tmp12047;
	wire signed [31:0] w_sys_tmp12048;
	wire signed [31:0] w_sys_tmp12052;
	wire signed [31:0] w_sys_tmp12053;
	wire signed [31:0] w_sys_tmp12057;
	wire signed [31:0] w_sys_tmp12058;
	wire signed [31:0] w_sys_tmp12062;
	wire signed [31:0] w_sys_tmp12063;
	wire signed [31:0] w_sys_tmp12067;
	wire signed [31:0] w_sys_tmp12068;
	wire signed [31:0] w_sys_tmp12072;
	wire signed [31:0] w_sys_tmp12073;
	wire signed [31:0] w_sys_tmp12077;
	wire signed [31:0] w_sys_tmp12078;
	wire signed [31:0] w_sys_tmp12082;
	wire signed [31:0] w_sys_tmp12083;
	wire signed [31:0] w_sys_tmp12087;
	wire signed [31:0] w_sys_tmp12088;
	wire signed [31:0] w_sys_tmp12092;
	wire signed [31:0] w_sys_tmp12093;
	wire signed [31:0] w_sys_tmp12097;
	wire signed [31:0] w_sys_tmp12098;
	wire signed [31:0] w_sys_tmp12102;
	wire signed [31:0] w_sys_tmp12103;
	wire signed [31:0] w_sys_tmp12107;
	wire signed [31:0] w_sys_tmp12108;
	wire signed [31:0] w_sys_tmp12112;
	wire signed [31:0] w_sys_tmp12113;
	wire signed [31:0] w_sys_tmp12117;
	wire signed [31:0] w_sys_tmp12118;
	wire signed [31:0] w_sys_tmp12122;
	wire signed [31:0] w_sys_tmp12123;
	wire signed [31:0] w_sys_tmp12127;
	wire signed [31:0] w_sys_tmp12128;
	wire signed [31:0] w_sys_tmp12132;
	wire signed [31:0] w_sys_tmp12133;
	wire signed [31:0] w_sys_tmp12137;
	wire signed [31:0] w_sys_tmp12138;
	wire signed [31:0] w_sys_tmp12142;
	wire signed [31:0] w_sys_tmp12143;
	wire signed [31:0] w_sys_tmp12147;
	wire signed [31:0] w_sys_tmp12148;
	wire signed [31:0] w_sys_tmp12152;
	wire signed [31:0] w_sys_tmp12153;
	wire signed [31:0] w_sys_tmp12157;
	wire signed [31:0] w_sys_tmp12158;
	wire signed [31:0] w_sys_tmp12162;
	wire signed [31:0] w_sys_tmp12163;
	wire signed [31:0] w_sys_tmp12167;
	wire signed [31:0] w_sys_tmp12168;
	wire signed [31:0] w_sys_tmp12172;
	wire signed [31:0] w_sys_tmp12173;
	wire signed [31:0] w_sys_tmp12177;
	wire signed [31:0] w_sys_tmp12178;
	wire signed [31:0] w_sys_tmp12182;
	wire signed [31:0] w_sys_tmp12183;
	wire signed [31:0] w_sys_tmp12187;
	wire signed [31:0] w_sys_tmp12188;
	wire signed [31:0] w_sys_tmp12192;
	wire signed [31:0] w_sys_tmp12193;
	wire signed [31:0] w_sys_tmp12197;
	wire signed [31:0] w_sys_tmp12198;
	wire signed [31:0] w_sys_tmp12202;
	wire signed [31:0] w_sys_tmp12203;
	wire signed [31:0] w_sys_tmp12207;
	wire signed [31:0] w_sys_tmp12208;
	wire signed [31:0] w_sys_tmp12212;
	wire signed [31:0] w_sys_tmp12213;
	wire signed [31:0] w_sys_tmp12217;
	wire signed [31:0] w_sys_tmp12218;
	wire signed [31:0] w_sys_tmp12222;
	wire signed [31:0] w_sys_tmp12223;
	wire signed [31:0] w_sys_tmp12227;
	wire signed [31:0] w_sys_tmp12228;
	wire signed [31:0] w_sys_tmp12232;
	wire signed [31:0] w_sys_tmp12233;
	wire signed [31:0] w_sys_tmp12237;
	wire signed [31:0] w_sys_tmp12238;
	wire signed [31:0] w_sys_tmp12242;
	wire signed [31:0] w_sys_tmp12243;
	wire signed [31:0] w_sys_tmp12247;
	wire signed [31:0] w_sys_tmp12248;
	wire signed [31:0] w_sys_tmp12252;
	wire signed [31:0] w_sys_tmp12253;
	wire signed [31:0] w_sys_tmp12257;
	wire signed [31:0] w_sys_tmp12258;
	wire signed [31:0] w_sys_tmp12262;
	wire signed [31:0] w_sys_tmp12263;
	wire signed [31:0] w_sys_tmp12267;
	wire signed [31:0] w_sys_tmp12268;
	wire signed [31:0] w_sys_tmp12272;
	wire signed [31:0] w_sys_tmp12273;
	wire signed [31:0] w_sys_tmp12277;
	wire signed [31:0] w_sys_tmp12278;
	wire signed [31:0] w_sys_tmp12282;
	wire signed [31:0] w_sys_tmp12283;
	wire signed [31:0] w_sys_tmp12287;
	wire signed [31:0] w_sys_tmp12288;
	wire signed [31:0] w_sys_tmp12292;
	wire signed [31:0] w_sys_tmp12293;
	wire signed [31:0] w_sys_tmp12297;
	wire signed [31:0] w_sys_tmp12298;
	wire signed [31:0] w_sys_tmp12302;
	wire signed [31:0] w_sys_tmp12303;
	wire signed [31:0] w_sys_tmp12307;
	wire signed [31:0] w_sys_tmp12308;
	wire signed [31:0] w_sys_tmp12312;
	wire signed [31:0] w_sys_tmp12313;
	wire signed [31:0] w_sys_tmp12317;
	wire signed [31:0] w_sys_tmp12318;
	wire signed [31:0] w_sys_tmp12322;
	wire signed [31:0] w_sys_tmp12323;
	wire signed [31:0] w_sys_tmp12327;
	wire signed [31:0] w_sys_tmp12328;
	wire signed [31:0] w_sys_tmp12332;
	wire signed [31:0] w_sys_tmp12333;
	wire signed [31:0] w_sys_tmp12337;
	wire signed [31:0] w_sys_tmp12338;
	wire signed [31:0] w_sys_tmp12342;
	wire signed [31:0] w_sys_tmp12343;
	wire signed [31:0] w_sys_tmp12347;
	wire signed [31:0] w_sys_tmp12348;
	wire signed [31:0] w_sys_tmp12352;
	wire signed [31:0] w_sys_tmp12353;
	wire signed [31:0] w_sys_tmp12357;
	wire signed [31:0] w_sys_tmp12358;
	wire signed [31:0] w_sys_tmp12362;
	wire signed [31:0] w_sys_tmp12363;
	wire signed [31:0] w_sys_tmp12367;
	wire signed [31:0] w_sys_tmp12368;
	wire signed [31:0] w_sys_tmp12372;
	wire signed [31:0] w_sys_tmp12373;
	wire signed [31:0] w_sys_tmp12377;
	wire signed [31:0] w_sys_tmp12378;
	wire signed [31:0] w_sys_tmp12382;
	wire signed [31:0] w_sys_tmp12383;
	wire signed [31:0] w_sys_tmp12387;
	wire signed [31:0] w_sys_tmp12388;
	wire signed [31:0] w_sys_tmp12392;
	wire signed [31:0] w_sys_tmp12393;
	wire signed [31:0] w_sys_tmp12397;
	wire signed [31:0] w_sys_tmp12398;
	wire signed [31:0] w_sys_tmp12402;
	wire signed [31:0] w_sys_tmp12403;
	wire signed [31:0] w_sys_tmp12407;
	wire signed [31:0] w_sys_tmp12408;
	wire signed [31:0] w_sys_tmp12412;
	wire signed [31:0] w_sys_tmp12413;
	wire signed [31:0] w_sys_tmp12417;
	wire signed [31:0] w_sys_tmp12418;
	wire signed [31:0] w_sys_tmp12422;
	wire signed [31:0] w_sys_tmp12423;
	wire signed [31:0] w_sys_tmp12427;
	wire signed [31:0] w_sys_tmp12428;
	wire signed [31:0] w_sys_tmp12432;
	wire signed [31:0] w_sys_tmp12433;
	wire signed [31:0] w_sys_tmp12437;
	wire signed [31:0] w_sys_tmp12438;
	wire signed [31:0] w_sys_tmp12442;
	wire signed [31:0] w_sys_tmp12443;
	wire signed [31:0] w_sys_tmp12447;
	wire signed [31:0] w_sys_tmp12448;
	wire signed [31:0] w_sys_tmp12452;
	wire signed [31:0] w_sys_tmp12453;
	wire signed [31:0] w_sys_tmp12457;
	wire signed [31:0] w_sys_tmp12458;
	wire signed [31:0] w_sys_tmp12462;
	wire signed [31:0] w_sys_tmp12463;
	wire signed [31:0] w_sys_tmp12467;
	wire signed [31:0] w_sys_tmp12468;
	wire signed [31:0] w_sys_tmp12472;
	wire signed [31:0] w_sys_tmp12473;
	wire signed [31:0] w_sys_tmp12477;
	wire signed [31:0] w_sys_tmp12478;
	wire signed [31:0] w_sys_tmp12482;
	wire signed [31:0] w_sys_tmp12483;
	wire signed [31:0] w_sys_tmp12487;
	wire signed [31:0] w_sys_tmp12488;
	wire signed [31:0] w_sys_tmp12492;
	wire signed [31:0] w_sys_tmp12493;
	wire signed [31:0] w_sys_tmp12497;
	wire signed [31:0] w_sys_tmp12498;
	wire signed [31:0] w_sys_tmp12502;
	wire signed [31:0] w_sys_tmp12503;
	wire signed [31:0] w_sys_tmp12507;
	wire signed [31:0] w_sys_tmp12508;
	wire signed [31:0] w_sys_tmp12512;
	wire signed [31:0] w_sys_tmp12513;
	wire signed [31:0] w_sys_tmp12517;
	wire signed [31:0] w_sys_tmp12518;
	wire signed [31:0] w_sys_tmp12522;
	wire signed [31:0] w_sys_tmp12523;
	wire signed [31:0] w_sys_tmp12527;
	wire signed [31:0] w_sys_tmp12528;
	wire signed [31:0] w_sys_tmp12532;
	wire signed [31:0] w_sys_tmp12533;
	wire signed [31:0] w_sys_tmp12537;
	wire signed [31:0] w_sys_tmp12538;
	wire signed [31:0] w_sys_tmp12542;
	wire signed [31:0] w_sys_tmp12543;
	wire signed [31:0] w_sys_tmp12547;
	wire signed [31:0] w_sys_tmp12548;
	wire signed [31:0] w_sys_tmp12552;
	wire signed [31:0] w_sys_tmp12553;
	wire signed [31:0] w_sys_tmp12557;
	wire signed [31:0] w_sys_tmp12558;
	wire signed [31:0] w_sys_tmp12562;
	wire signed [31:0] w_sys_tmp12563;
	wire signed [31:0] w_sys_tmp12567;
	wire signed [31:0] w_sys_tmp12568;
	wire signed [31:0] w_sys_tmp12572;
	wire signed [31:0] w_sys_tmp12573;
	wire signed [31:0] w_sys_tmp12577;
	wire signed [31:0] w_sys_tmp12578;
	wire signed [31:0] w_sys_tmp12582;
	wire signed [31:0] w_sys_tmp12583;
	wire signed [31:0] w_sys_tmp12587;
	wire signed [31:0] w_sys_tmp12588;
	wire signed [31:0] w_sys_tmp12592;
	wire signed [31:0] w_sys_tmp12593;
	wire signed [31:0] w_sys_tmp12597;
	wire signed [31:0] w_sys_tmp12598;
	wire signed [31:0] w_sys_tmp12602;
	wire signed [31:0] w_sys_tmp12603;
	wire signed [31:0] w_sys_tmp12607;
	wire signed [31:0] w_sys_tmp12608;
	wire signed [31:0] w_sys_tmp12612;
	wire signed [31:0] w_sys_tmp12613;
	wire signed [31:0] w_sys_tmp12617;
	wire signed [31:0] w_sys_tmp12618;
	wire signed [31:0] w_sys_tmp12622;
	wire signed [31:0] w_sys_tmp12623;
	wire signed [31:0] w_sys_tmp12627;
	wire signed [31:0] w_sys_tmp12628;
	wire signed [31:0] w_sys_tmp12632;
	wire signed [31:0] w_sys_tmp12633;
	wire signed [31:0] w_sys_tmp12637;
	wire signed [31:0] w_sys_tmp12638;
	wire signed [31:0] w_sys_tmp12642;
	wire signed [31:0] w_sys_tmp12643;
	wire signed [31:0] w_sys_tmp12647;
	wire signed [31:0] w_sys_tmp12648;
	wire signed [31:0] w_sys_tmp12652;
	wire signed [31:0] w_sys_tmp12653;
	wire signed [31:0] w_sys_tmp12657;
	wire signed [31:0] w_sys_tmp12658;
	wire signed [31:0] w_sys_tmp12662;
	wire signed [31:0] w_sys_tmp12663;
	wire signed [31:0] w_sys_tmp12667;
	wire signed [31:0] w_sys_tmp12668;
	wire signed [31:0] w_sys_tmp12672;
	wire signed [31:0] w_sys_tmp12673;
	wire signed [31:0] w_sys_tmp12677;
	wire signed [31:0] w_sys_tmp12678;
	wire signed [31:0] w_sys_tmp12682;
	wire signed [31:0] w_sys_tmp12683;
	wire signed [31:0] w_sys_tmp12687;
	wire signed [31:0] w_sys_tmp12688;
	wire signed [31:0] w_sys_tmp12692;
	wire signed [31:0] w_sys_tmp12693;
	wire signed [31:0] w_sys_tmp12697;
	wire signed [31:0] w_sys_tmp12698;
	wire signed [31:0] w_sys_tmp12702;
	wire signed [31:0] w_sys_tmp12703;
	wire signed [31:0] w_sys_tmp12707;
	wire signed [31:0] w_sys_tmp12708;
	wire signed [31:0] w_sys_tmp12712;
	wire signed [31:0] w_sys_tmp12713;
	wire signed [31:0] w_sys_tmp12717;
	wire signed [31:0] w_sys_tmp12718;
	wire signed [31:0] w_sys_tmp12722;
	wire signed [31:0] w_sys_tmp12723;
	wire signed [31:0] w_sys_tmp12727;
	wire signed [31:0] w_sys_tmp12728;
	wire signed [31:0] w_sys_tmp12732;
	wire signed [31:0] w_sys_tmp12733;
	wire signed [31:0] w_sys_tmp12737;
	wire signed [31:0] w_sys_tmp12738;
	wire signed [31:0] w_sys_tmp12742;
	wire signed [31:0] w_sys_tmp12743;
	wire signed [31:0] w_sys_tmp12747;
	wire signed [31:0] w_sys_tmp12748;
	wire signed [31:0] w_sys_tmp12752;
	wire signed [31:0] w_sys_tmp12753;
	wire signed [31:0] w_sys_tmp12757;
	wire signed [31:0] w_sys_tmp12758;
	wire signed [31:0] w_sys_tmp12762;
	wire signed [31:0] w_sys_tmp12763;
	wire signed [31:0] w_sys_tmp12767;
	wire signed [31:0] w_sys_tmp12768;
	wire signed [31:0] w_sys_tmp12772;
	wire signed [31:0] w_sys_tmp12773;
	wire signed [31:0] w_sys_tmp12777;
	wire signed [31:0] w_sys_tmp12778;
	wire signed [31:0] w_sys_tmp12782;
	wire signed [31:0] w_sys_tmp12783;
	wire signed [31:0] w_sys_tmp12787;
	wire signed [31:0] w_sys_tmp12788;
	wire signed [31:0] w_sys_tmp12792;
	wire signed [31:0] w_sys_tmp12793;
	wire signed [31:0] w_sys_tmp12797;
	wire signed [31:0] w_sys_tmp12798;
	wire signed [31:0] w_sys_tmp12802;
	wire signed [31:0] w_sys_tmp12803;
	wire signed [31:0] w_sys_tmp12807;
	wire signed [31:0] w_sys_tmp12808;
	wire signed [31:0] w_sys_tmp12812;
	wire signed [31:0] w_sys_tmp12813;
	wire signed [31:0] w_sys_tmp12817;
	wire signed [31:0] w_sys_tmp12818;
	wire signed [31:0] w_sys_tmp12822;
	wire signed [31:0] w_sys_tmp12823;
	wire signed [31:0] w_sys_tmp12827;
	wire signed [31:0] w_sys_tmp12828;
	wire signed [31:0] w_sys_tmp12832;
	wire signed [31:0] w_sys_tmp12833;
	wire signed [31:0] w_sys_tmp12837;
	wire signed [31:0] w_sys_tmp12838;
	wire signed [31:0] w_sys_tmp12842;
	wire signed [31:0] w_sys_tmp12843;
	wire signed [31:0] w_sys_tmp12847;
	wire signed [31:0] w_sys_tmp12848;
	wire signed [31:0] w_sys_tmp12852;
	wire signed [31:0] w_sys_tmp12853;
	wire signed [31:0] w_sys_tmp12857;
	wire signed [31:0] w_sys_tmp12858;
	wire signed [31:0] w_sys_tmp12862;
	wire signed [31:0] w_sys_tmp12863;
	wire signed [31:0] w_sys_tmp12867;
	wire signed [31:0] w_sys_tmp12868;
	wire signed [31:0] w_sys_tmp12872;
	wire signed [31:0] w_sys_tmp12873;
	wire signed [31:0] w_sys_tmp12877;
	wire signed [31:0] w_sys_tmp12878;
	wire signed [31:0] w_sys_tmp12882;
	wire signed [31:0] w_sys_tmp12883;
	wire signed [31:0] w_sys_tmp12887;
	wire signed [31:0] w_sys_tmp12888;
	wire signed [31:0] w_sys_tmp12892;
	wire signed [31:0] w_sys_tmp12893;
	wire signed [31:0] w_sys_tmp12897;
	wire signed [31:0] w_sys_tmp12898;
	wire signed [31:0] w_sys_tmp12902;
	wire signed [31:0] w_sys_tmp12903;
	wire signed [31:0] w_sys_tmp12907;
	wire signed [31:0] w_sys_tmp12908;
	wire signed [31:0] w_sys_tmp12912;
	wire signed [31:0] w_sys_tmp12913;
	wire signed [31:0] w_sys_tmp12917;
	wire signed [31:0] w_sys_tmp12918;
	wire signed [31:0] w_sys_tmp12922;
	wire signed [31:0] w_sys_tmp12923;
	wire signed [31:0] w_sys_tmp12927;
	wire signed [31:0] w_sys_tmp12928;
	wire signed [31:0] w_sys_tmp12932;
	wire signed [31:0] w_sys_tmp12933;
	wire signed [31:0] w_sys_tmp12937;
	wire signed [31:0] w_sys_tmp12938;
	wire signed [31:0] w_sys_tmp12942;
	wire signed [31:0] w_sys_tmp12943;
	wire signed [31:0] w_sys_tmp12947;
	wire signed [31:0] w_sys_tmp12948;
	wire signed [31:0] w_sys_tmp12951;
	wire signed [31:0] w_sys_tmp12952;
	wire               w_sys_tmp12953;
	wire               w_sys_tmp12954;
	wire signed [31:0] w_sys_tmp12955;
	wire signed [31:0] w_sys_tmp12958;
	wire signed [31:0] w_sys_tmp12959;
	wire        [31:0] w_sys_tmp12960;
	wire signed [31:0] w_sys_tmp12964;
	wire signed [31:0] w_sys_tmp12965;
	wire signed [31:0] w_sys_tmp12970;
	wire signed [31:0] w_sys_tmp12971;
	wire signed [31:0] w_sys_tmp12976;
	wire signed [31:0] w_sys_tmp12977;
	wire signed [31:0] w_sys_tmp12982;
	wire signed [31:0] w_sys_tmp12983;
	wire signed [31:0] w_sys_tmp12988;
	wire signed [31:0] w_sys_tmp12989;
	wire signed [31:0] w_sys_tmp12994;
	wire signed [31:0] w_sys_tmp12995;
	wire signed [31:0] w_sys_tmp13000;
	wire signed [31:0] w_sys_tmp13001;
	wire signed [31:0] w_sys_tmp13006;
	wire signed [31:0] w_sys_tmp13007;
	wire signed [31:0] w_sys_tmp13012;
	wire signed [31:0] w_sys_tmp13013;
	wire signed [31:0] w_sys_tmp13018;
	wire signed [31:0] w_sys_tmp13019;
	wire signed [31:0] w_sys_tmp13024;
	wire signed [31:0] w_sys_tmp13025;
	wire signed [31:0] w_sys_tmp13030;
	wire signed [31:0] w_sys_tmp13031;
	wire signed [31:0] w_sys_tmp13036;
	wire signed [31:0] w_sys_tmp13037;
	wire signed [31:0] w_sys_tmp13042;
	wire signed [31:0] w_sys_tmp13043;
	wire signed [31:0] w_sys_tmp13048;
	wire signed [31:0] w_sys_tmp13049;
	wire signed [31:0] w_sys_tmp13054;
	wire signed [31:0] w_sys_tmp13055;
	wire signed [31:0] w_sys_tmp13060;
	wire signed [31:0] w_sys_tmp13061;
	wire signed [31:0] w_sys_tmp13066;
	wire signed [31:0] w_sys_tmp13067;
	wire signed [31:0] w_sys_tmp13072;
	wire signed [31:0] w_sys_tmp13073;
	wire signed [31:0] w_sys_tmp13078;
	wire signed [31:0] w_sys_tmp13079;
	wire signed [31:0] w_sys_tmp13083;
	wire signed [31:0] w_sys_tmp13084;
	wire signed [31:0] w_sys_tmp13088;
	wire signed [31:0] w_sys_tmp13089;
	wire signed [31:0] w_sys_tmp13093;
	wire signed [31:0] w_sys_tmp13094;
	wire signed [31:0] w_sys_tmp13098;
	wire signed [31:0] w_sys_tmp13099;
	wire signed [31:0] w_sys_tmp13103;
	wire signed [31:0] w_sys_tmp13104;
	wire signed [31:0] w_sys_tmp13108;
	wire signed [31:0] w_sys_tmp13109;
	wire signed [31:0] w_sys_tmp13113;
	wire signed [31:0] w_sys_tmp13114;
	wire signed [31:0] w_sys_tmp13118;
	wire signed [31:0] w_sys_tmp13119;
	wire signed [31:0] w_sys_tmp13123;
	wire signed [31:0] w_sys_tmp13124;
	wire signed [31:0] w_sys_tmp13128;
	wire signed [31:0] w_sys_tmp13129;
	wire signed [31:0] w_sys_tmp13133;
	wire signed [31:0] w_sys_tmp13134;
	wire signed [31:0] w_sys_tmp13138;
	wire signed [31:0] w_sys_tmp13139;
	wire signed [31:0] w_sys_tmp13143;
	wire signed [31:0] w_sys_tmp13144;
	wire signed [31:0] w_sys_tmp13148;
	wire signed [31:0] w_sys_tmp13149;
	wire signed [31:0] w_sys_tmp13153;
	wire signed [31:0] w_sys_tmp13154;
	wire signed [31:0] w_sys_tmp13158;
	wire signed [31:0] w_sys_tmp13159;
	wire signed [31:0] w_sys_tmp13163;
	wire signed [31:0] w_sys_tmp13164;
	wire signed [31:0] w_sys_tmp13168;
	wire signed [31:0] w_sys_tmp13169;
	wire signed [31:0] w_sys_tmp13173;
	wire signed [31:0] w_sys_tmp13174;
	wire signed [31:0] w_sys_tmp13178;
	wire signed [31:0] w_sys_tmp13179;
	wire signed [31:0] w_sys_tmp13183;
	wire signed [31:0] w_sys_tmp13184;
	wire signed [31:0] w_sys_tmp13188;
	wire signed [31:0] w_sys_tmp13189;
	wire signed [31:0] w_sys_tmp13193;
	wire signed [31:0] w_sys_tmp13194;
	wire signed [31:0] w_sys_tmp13198;
	wire signed [31:0] w_sys_tmp13199;
	wire signed [31:0] w_sys_tmp13203;
	wire signed [31:0] w_sys_tmp13204;
	wire signed [31:0] w_sys_tmp13208;
	wire signed [31:0] w_sys_tmp13209;
	wire signed [31:0] w_sys_tmp13213;
	wire signed [31:0] w_sys_tmp13214;
	wire signed [31:0] w_sys_tmp13218;
	wire signed [31:0] w_sys_tmp13219;
	wire signed [31:0] w_sys_tmp13223;
	wire signed [31:0] w_sys_tmp13224;
	wire signed [31:0] w_sys_tmp13228;
	wire signed [31:0] w_sys_tmp13229;
	wire signed [31:0] w_sys_tmp13233;
	wire signed [31:0] w_sys_tmp13234;
	wire signed [31:0] w_sys_tmp13238;
	wire signed [31:0] w_sys_tmp13239;
	wire signed [31:0] w_sys_tmp13243;
	wire signed [31:0] w_sys_tmp13244;
	wire signed [31:0] w_sys_tmp13248;
	wire signed [31:0] w_sys_tmp13249;
	wire signed [31:0] w_sys_tmp13253;
	wire signed [31:0] w_sys_tmp13254;
	wire signed [31:0] w_sys_tmp13258;
	wire signed [31:0] w_sys_tmp13259;
	wire signed [31:0] w_sys_tmp13263;
	wire signed [31:0] w_sys_tmp13264;
	wire signed [31:0] w_sys_tmp13268;
	wire signed [31:0] w_sys_tmp13269;
	wire signed [31:0] w_sys_tmp13273;
	wire signed [31:0] w_sys_tmp13274;
	wire signed [31:0] w_sys_tmp13278;
	wire signed [31:0] w_sys_tmp13279;
	wire signed [31:0] w_sys_tmp13283;
	wire signed [31:0] w_sys_tmp13284;
	wire signed [31:0] w_sys_tmp13288;
	wire signed [31:0] w_sys_tmp13289;
	wire signed [31:0] w_sys_tmp13293;
	wire signed [31:0] w_sys_tmp13294;
	wire signed [31:0] w_sys_tmp13298;
	wire signed [31:0] w_sys_tmp13299;
	wire signed [31:0] w_sys_tmp13303;
	wire signed [31:0] w_sys_tmp13304;
	wire signed [31:0] w_sys_tmp13308;
	wire signed [31:0] w_sys_tmp13309;
	wire signed [31:0] w_sys_tmp13313;
	wire signed [31:0] w_sys_tmp13314;
	wire signed [31:0] w_sys_tmp13318;
	wire signed [31:0] w_sys_tmp13319;
	wire signed [31:0] w_sys_tmp13323;
	wire signed [31:0] w_sys_tmp13324;
	wire signed [31:0] w_sys_tmp13328;
	wire signed [31:0] w_sys_tmp13329;
	wire signed [31:0] w_sys_tmp13333;
	wire signed [31:0] w_sys_tmp13334;
	wire signed [31:0] w_sys_tmp13338;
	wire signed [31:0] w_sys_tmp13339;
	wire signed [31:0] w_sys_tmp13343;
	wire signed [31:0] w_sys_tmp13344;
	wire signed [31:0] w_sys_tmp13348;
	wire signed [31:0] w_sys_tmp13349;
	wire signed [31:0] w_sys_tmp13353;
	wire signed [31:0] w_sys_tmp13354;
	wire signed [31:0] w_sys_tmp13358;
	wire signed [31:0] w_sys_tmp13359;
	wire signed [31:0] w_sys_tmp13363;
	wire signed [31:0] w_sys_tmp13364;
	wire signed [31:0] w_sys_tmp13368;
	wire signed [31:0] w_sys_tmp13369;
	wire signed [31:0] w_sys_tmp13373;
	wire signed [31:0] w_sys_tmp13374;
	wire signed [31:0] w_sys_tmp13378;
	wire signed [31:0] w_sys_tmp13379;
	wire signed [31:0] w_sys_tmp13383;
	wire signed [31:0] w_sys_tmp13384;
	wire signed [31:0] w_sys_tmp13388;
	wire signed [31:0] w_sys_tmp13389;
	wire signed [31:0] w_sys_tmp13393;
	wire signed [31:0] w_sys_tmp13394;
	wire signed [31:0] w_sys_tmp13398;
	wire signed [31:0] w_sys_tmp13399;
	wire signed [31:0] w_sys_tmp13403;
	wire signed [31:0] w_sys_tmp13404;
	wire signed [31:0] w_sys_tmp13408;
	wire signed [31:0] w_sys_tmp13409;
	wire signed [31:0] w_sys_tmp13413;
	wire signed [31:0] w_sys_tmp13414;
	wire signed [31:0] w_sys_tmp13418;
	wire signed [31:0] w_sys_tmp13419;
	wire signed [31:0] w_sys_tmp13423;
	wire signed [31:0] w_sys_tmp13424;
	wire signed [31:0] w_sys_tmp13428;
	wire signed [31:0] w_sys_tmp13429;
	wire signed [31:0] w_sys_tmp13433;
	wire signed [31:0] w_sys_tmp13434;
	wire signed [31:0] w_sys_tmp13438;
	wire signed [31:0] w_sys_tmp13439;
	wire signed [31:0] w_sys_tmp13443;
	wire signed [31:0] w_sys_tmp13444;
	wire signed [31:0] w_sys_tmp13448;
	wire signed [31:0] w_sys_tmp13449;
	wire signed [31:0] w_sys_tmp13453;
	wire signed [31:0] w_sys_tmp13454;
	wire signed [31:0] w_sys_tmp13458;
	wire signed [31:0] w_sys_tmp13459;
	wire signed [31:0] w_sys_tmp13463;
	wire signed [31:0] w_sys_tmp13464;
	wire signed [31:0] w_sys_tmp13468;
	wire signed [31:0] w_sys_tmp13469;
	wire signed [31:0] w_sys_tmp13472;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 5'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 9'h1);
	assign w_fld_T_0_addr_0 = 14'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 14'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 14'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_fld_V_3_addr_0 = 14'sh0;
	assign w_fld_V_3_datain_0 = 32'h0;
	assign w_fld_V_3_r_w_0 = 1'h0;
	assign w_fld_V_3_ce_0 = w_sys_ce;
	assign w_fld_V_3_ce_1 = w_sys_ce;
	assign w_sub19_T_addr = ( (|r_sys_processing_methodID) ? r_sub19_T_addr : 14'sh0 ) ;
	assign w_sub19_T_datain = ( (|r_sys_processing_methodID) ? r_sub19_T_datain : 32'h0 ) ;
	assign w_sub19_T_r_w = ( (|r_sys_processing_methodID) ? r_sub19_T_r_w : 1'h0 ) ;
	assign w_sub19_V_addr = ( (|r_sys_processing_methodID) ? r_sub19_V_addr : 14'sh0 ) ;
	assign w_sub19_V_datain = ( (|r_sys_processing_methodID) ? r_sub19_V_datain : 32'h0 ) ;
	assign w_sub19_V_r_w = ( (|r_sys_processing_methodID) ? r_sub19_V_r_w : 1'h0 ) ;
	assign w_sub19_U_addr = ( (|r_sys_processing_methodID) ? r_sub19_U_addr : 14'sh0 ) ;
	assign w_sub19_U_datain = ( (|r_sys_processing_methodID) ? r_sub19_U_datain : 32'h0 ) ;
	assign w_sub19_U_r_w = ( (|r_sys_processing_methodID) ? r_sub19_U_r_w : 1'h0 ) ;
	assign w_sub19_result_addr = ( (|r_sys_processing_methodID) ? r_sub19_result_addr : 14'sh0 ) ;
	assign w_sub19_result_datain = ( (|r_sys_processing_methodID) ? r_sub19_result_datain : 32'h0 ) ;
	assign w_sub19_result_r_w = ( (|r_sys_processing_methodID) ? r_sub19_result_r_w : 1'h0 ) ;
	assign w_sub09_T_addr = ( (|r_sys_processing_methodID) ? r_sub09_T_addr : 14'sh0 ) ;
	assign w_sub09_T_datain = ( (|r_sys_processing_methodID) ? r_sub09_T_datain : 32'h0 ) ;
	assign w_sub09_T_r_w = ( (|r_sys_processing_methodID) ? r_sub09_T_r_w : 1'h0 ) ;
	assign w_sub09_V_addr = ( (|r_sys_processing_methodID) ? r_sub09_V_addr : 14'sh0 ) ;
	assign w_sub09_V_datain = ( (|r_sys_processing_methodID) ? r_sub09_V_datain : 32'h0 ) ;
	assign w_sub09_V_r_w = ( (|r_sys_processing_methodID) ? r_sub09_V_r_w : 1'h0 ) ;
	assign w_sub09_U_addr = ( (|r_sys_processing_methodID) ? r_sub09_U_addr : 14'sh0 ) ;
	assign w_sub09_U_datain = ( (|r_sys_processing_methodID) ? r_sub09_U_datain : 32'h0 ) ;
	assign w_sub09_U_r_w = ( (|r_sys_processing_methodID) ? r_sub09_U_r_w : 1'h0 ) ;
	assign w_sub09_result_addr = ( (|r_sys_processing_methodID) ? r_sub09_result_addr : 14'sh0 ) ;
	assign w_sub09_result_datain = ( (|r_sys_processing_methodID) ? r_sub09_result_datain : 32'h0 ) ;
	assign w_sub09_result_r_w = ( (|r_sys_processing_methodID) ? r_sub09_result_r_w : 1'h0 ) ;
	assign w_sub08_T_addr = ( (|r_sys_processing_methodID) ? r_sub08_T_addr : 14'sh0 ) ;
	assign w_sub08_T_datain = ( (|r_sys_processing_methodID) ? r_sub08_T_datain : 32'h0 ) ;
	assign w_sub08_T_r_w = ( (|r_sys_processing_methodID) ? r_sub08_T_r_w : 1'h0 ) ;
	assign w_sub08_V_addr = ( (|r_sys_processing_methodID) ? r_sub08_V_addr : 14'sh0 ) ;
	assign w_sub08_V_datain = ( (|r_sys_processing_methodID) ? r_sub08_V_datain : 32'h0 ) ;
	assign w_sub08_V_r_w = ( (|r_sys_processing_methodID) ? r_sub08_V_r_w : 1'h0 ) ;
	assign w_sub08_U_addr = ( (|r_sys_processing_methodID) ? r_sub08_U_addr : 14'sh0 ) ;
	assign w_sub08_U_datain = ( (|r_sys_processing_methodID) ? r_sub08_U_datain : 32'h0 ) ;
	assign w_sub08_U_r_w = ( (|r_sys_processing_methodID) ? r_sub08_U_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 14'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub24_T_addr = ( (|r_sys_processing_methodID) ? r_sub24_T_addr : 14'sh0 ) ;
	assign w_sub24_T_datain = ( (|r_sys_processing_methodID) ? r_sub24_T_datain : 32'h0 ) ;
	assign w_sub24_T_r_w = ( (|r_sys_processing_methodID) ? r_sub24_T_r_w : 1'h0 ) ;
	assign w_sub24_V_addr = ( (|r_sys_processing_methodID) ? r_sub24_V_addr : 14'sh0 ) ;
	assign w_sub24_V_datain = ( (|r_sys_processing_methodID) ? r_sub24_V_datain : 32'h0 ) ;
	assign w_sub24_V_r_w = ( (|r_sys_processing_methodID) ? r_sub24_V_r_w : 1'h0 ) ;
	assign w_sub24_U_addr = ( (|r_sys_processing_methodID) ? r_sub24_U_addr : 14'sh0 ) ;
	assign w_sub24_U_datain = ( (|r_sys_processing_methodID) ? r_sub24_U_datain : 32'h0 ) ;
	assign w_sub24_U_r_w = ( (|r_sys_processing_methodID) ? r_sub24_U_r_w : 1'h0 ) ;
	assign w_sub24_result_addr = ( (|r_sys_processing_methodID) ? r_sub24_result_addr : 14'sh0 ) ;
	assign w_sub24_result_datain = ( (|r_sys_processing_methodID) ? r_sub24_result_datain : 32'h0 ) ;
	assign w_sub24_result_r_w = ( (|r_sys_processing_methodID) ? r_sub24_result_r_w : 1'h0 ) ;
	assign w_sub22_T_addr = ( (|r_sys_processing_methodID) ? r_sub22_T_addr : 14'sh0 ) ;
	assign w_sub22_T_datain = ( (|r_sys_processing_methodID) ? r_sub22_T_datain : 32'h0 ) ;
	assign w_sub22_T_r_w = ( (|r_sys_processing_methodID) ? r_sub22_T_r_w : 1'h0 ) ;
	assign w_sub22_V_addr = ( (|r_sys_processing_methodID) ? r_sub22_V_addr : 14'sh0 ) ;
	assign w_sub22_V_datain = ( (|r_sys_processing_methodID) ? r_sub22_V_datain : 32'h0 ) ;
	assign w_sub22_V_r_w = ( (|r_sys_processing_methodID) ? r_sub22_V_r_w : 1'h0 ) ;
	assign w_sub22_U_addr = ( (|r_sys_processing_methodID) ? r_sub22_U_addr : 14'sh0 ) ;
	assign w_sub22_U_datain = ( (|r_sys_processing_methodID) ? r_sub22_U_datain : 32'h0 ) ;
	assign w_sub22_U_r_w = ( (|r_sys_processing_methodID) ? r_sub22_U_r_w : 1'h0 ) ;
	assign w_sub22_result_addr = ( (|r_sys_processing_methodID) ? r_sub22_result_addr : 14'sh0 ) ;
	assign w_sub22_result_datain = ( (|r_sys_processing_methodID) ? r_sub22_result_datain : 32'h0 ) ;
	assign w_sub22_result_r_w = ( (|r_sys_processing_methodID) ? r_sub22_result_r_w : 1'h0 ) ;
	assign w_sub23_T_addr = ( (|r_sys_processing_methodID) ? r_sub23_T_addr : 14'sh0 ) ;
	assign w_sub23_T_datain = ( (|r_sys_processing_methodID) ? r_sub23_T_datain : 32'h0 ) ;
	assign w_sub23_T_r_w = ( (|r_sys_processing_methodID) ? r_sub23_T_r_w : 1'h0 ) ;
	assign w_sub23_V_addr = ( (|r_sys_processing_methodID) ? r_sub23_V_addr : 14'sh0 ) ;
	assign w_sub23_V_datain = ( (|r_sys_processing_methodID) ? r_sub23_V_datain : 32'h0 ) ;
	assign w_sub23_V_r_w = ( (|r_sys_processing_methodID) ? r_sub23_V_r_w : 1'h0 ) ;
	assign w_sub23_U_addr = ( (|r_sys_processing_methodID) ? r_sub23_U_addr : 14'sh0 ) ;
	assign w_sub23_U_datain = ( (|r_sys_processing_methodID) ? r_sub23_U_datain : 32'h0 ) ;
	assign w_sub23_U_r_w = ( (|r_sys_processing_methodID) ? r_sub23_U_r_w : 1'h0 ) ;
	assign w_sub23_result_addr = ( (|r_sys_processing_methodID) ? r_sub23_result_addr : 14'sh0 ) ;
	assign w_sub23_result_datain = ( (|r_sys_processing_methodID) ? r_sub23_result_datain : 32'h0 ) ;
	assign w_sub23_result_r_w = ( (|r_sys_processing_methodID) ? r_sub23_result_r_w : 1'h0 ) ;
	assign w_sub12_T_addr = ( (|r_sys_processing_methodID) ? r_sub12_T_addr : 14'sh0 ) ;
	assign w_sub12_T_datain = ( (|r_sys_processing_methodID) ? r_sub12_T_datain : 32'h0 ) ;
	assign w_sub12_T_r_w = ( (|r_sys_processing_methodID) ? r_sub12_T_r_w : 1'h0 ) ;
	assign w_sub12_V_addr = ( (|r_sys_processing_methodID) ? r_sub12_V_addr : 14'sh0 ) ;
	assign w_sub12_V_datain = ( (|r_sys_processing_methodID) ? r_sub12_V_datain : 32'h0 ) ;
	assign w_sub12_V_r_w = ( (|r_sys_processing_methodID) ? r_sub12_V_r_w : 1'h0 ) ;
	assign w_sub12_U_addr = ( (|r_sys_processing_methodID) ? r_sub12_U_addr : 14'sh0 ) ;
	assign w_sub12_U_datain = ( (|r_sys_processing_methodID) ? r_sub12_U_datain : 32'h0 ) ;
	assign w_sub12_U_r_w = ( (|r_sys_processing_methodID) ? r_sub12_U_r_w : 1'h0 ) ;
	assign w_sub12_result_addr = ( (|r_sys_processing_methodID) ? r_sub12_result_addr : 14'sh0 ) ;
	assign w_sub12_result_datain = ( (|r_sys_processing_methodID) ? r_sub12_result_datain : 32'h0 ) ;
	assign w_sub12_result_r_w = ( (|r_sys_processing_methodID) ? r_sub12_result_r_w : 1'h0 ) ;
	assign w_sub03_T_addr = ( (|r_sys_processing_methodID) ? r_sub03_T_addr : 14'sh0 ) ;
	assign w_sub03_T_datain = ( (|r_sys_processing_methodID) ? r_sub03_T_datain : 32'h0 ) ;
	assign w_sub03_T_r_w = ( (|r_sys_processing_methodID) ? r_sub03_T_r_w : 1'h0 ) ;
	assign w_sub03_V_addr = ( (|r_sys_processing_methodID) ? r_sub03_V_addr : 14'sh0 ) ;
	assign w_sub03_V_datain = ( (|r_sys_processing_methodID) ? r_sub03_V_datain : 32'h0 ) ;
	assign w_sub03_V_r_w = ( (|r_sys_processing_methodID) ? r_sub03_V_r_w : 1'h0 ) ;
	assign w_sub03_U_addr = ( (|r_sys_processing_methodID) ? r_sub03_U_addr : 14'sh0 ) ;
	assign w_sub03_U_datain = ( (|r_sys_processing_methodID) ? r_sub03_U_datain : 32'h0 ) ;
	assign w_sub03_U_r_w = ( (|r_sys_processing_methodID) ? r_sub03_U_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 14'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_T_addr = ( (|r_sys_processing_methodID) ? r_sub02_T_addr : 14'sh0 ) ;
	assign w_sub02_T_datain = ( (|r_sys_processing_methodID) ? r_sub02_T_datain : 32'h0 ) ;
	assign w_sub02_T_r_w = ( (|r_sys_processing_methodID) ? r_sub02_T_r_w : 1'h0 ) ;
	assign w_sub02_V_addr = ( (|r_sys_processing_methodID) ? r_sub02_V_addr : 14'sh0 ) ;
	assign w_sub02_V_datain = ( (|r_sys_processing_methodID) ? r_sub02_V_datain : 32'h0 ) ;
	assign w_sub02_V_r_w = ( (|r_sys_processing_methodID) ? r_sub02_V_r_w : 1'h0 ) ;
	assign w_sub02_U_addr = ( (|r_sys_processing_methodID) ? r_sub02_U_addr : 14'sh0 ) ;
	assign w_sub02_U_datain = ( (|r_sys_processing_methodID) ? r_sub02_U_datain : 32'h0 ) ;
	assign w_sub02_U_r_w = ( (|r_sys_processing_methodID) ? r_sub02_U_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 14'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub11_T_addr = ( (|r_sys_processing_methodID) ? r_sub11_T_addr : 14'sh0 ) ;
	assign w_sub11_T_datain = ( (|r_sys_processing_methodID) ? r_sub11_T_datain : 32'h0 ) ;
	assign w_sub11_T_r_w = ( (|r_sys_processing_methodID) ? r_sub11_T_r_w : 1'h0 ) ;
	assign w_sub11_V_addr = ( (|r_sys_processing_methodID) ? r_sub11_V_addr : 14'sh0 ) ;
	assign w_sub11_V_datain = ( (|r_sys_processing_methodID) ? r_sub11_V_datain : 32'h0 ) ;
	assign w_sub11_V_r_w = ( (|r_sys_processing_methodID) ? r_sub11_V_r_w : 1'h0 ) ;
	assign w_sub11_U_addr = ( (|r_sys_processing_methodID) ? r_sub11_U_addr : 14'sh0 ) ;
	assign w_sub11_U_datain = ( (|r_sys_processing_methodID) ? r_sub11_U_datain : 32'h0 ) ;
	assign w_sub11_U_r_w = ( (|r_sys_processing_methodID) ? r_sub11_U_r_w : 1'h0 ) ;
	assign w_sub11_result_addr = ( (|r_sys_processing_methodID) ? r_sub11_result_addr : 14'sh0 ) ;
	assign w_sub11_result_datain = ( (|r_sys_processing_methodID) ? r_sub11_result_datain : 32'h0 ) ;
	assign w_sub11_result_r_w = ( (|r_sys_processing_methodID) ? r_sub11_result_r_w : 1'h0 ) ;
	assign w_sub14_T_addr = ( (|r_sys_processing_methodID) ? r_sub14_T_addr : 14'sh0 ) ;
	assign w_sub14_T_datain = ( (|r_sys_processing_methodID) ? r_sub14_T_datain : 32'h0 ) ;
	assign w_sub14_T_r_w = ( (|r_sys_processing_methodID) ? r_sub14_T_r_w : 1'h0 ) ;
	assign w_sub14_V_addr = ( (|r_sys_processing_methodID) ? r_sub14_V_addr : 14'sh0 ) ;
	assign w_sub14_V_datain = ( (|r_sys_processing_methodID) ? r_sub14_V_datain : 32'h0 ) ;
	assign w_sub14_V_r_w = ( (|r_sys_processing_methodID) ? r_sub14_V_r_w : 1'h0 ) ;
	assign w_sub14_U_addr = ( (|r_sys_processing_methodID) ? r_sub14_U_addr : 14'sh0 ) ;
	assign w_sub14_U_datain = ( (|r_sys_processing_methodID) ? r_sub14_U_datain : 32'h0 ) ;
	assign w_sub14_U_r_w = ( (|r_sys_processing_methodID) ? r_sub14_U_r_w : 1'h0 ) ;
	assign w_sub14_result_addr = ( (|r_sys_processing_methodID) ? r_sub14_result_addr : 14'sh0 ) ;
	assign w_sub14_result_datain = ( (|r_sys_processing_methodID) ? r_sub14_result_datain : 32'h0 ) ;
	assign w_sub14_result_r_w = ( (|r_sys_processing_methodID) ? r_sub14_result_r_w : 1'h0 ) ;
	assign w_sub01_T_addr = ( (|r_sys_processing_methodID) ? r_sub01_T_addr : 14'sh0 ) ;
	assign w_sub01_T_datain = ( (|r_sys_processing_methodID) ? r_sub01_T_datain : 32'h0 ) ;
	assign w_sub01_T_r_w = ( (|r_sys_processing_methodID) ? r_sub01_T_r_w : 1'h0 ) ;
	assign w_sub01_V_addr = ( (|r_sys_processing_methodID) ? r_sub01_V_addr : 14'sh0 ) ;
	assign w_sub01_V_datain = ( (|r_sys_processing_methodID) ? r_sub01_V_datain : 32'h0 ) ;
	assign w_sub01_V_r_w = ( (|r_sys_processing_methodID) ? r_sub01_V_r_w : 1'h0 ) ;
	assign w_sub01_U_addr = ( (|r_sys_processing_methodID) ? r_sub01_U_addr : 14'sh0 ) ;
	assign w_sub01_U_datain = ( (|r_sys_processing_methodID) ? r_sub01_U_datain : 32'h0 ) ;
	assign w_sub01_U_r_w = ( (|r_sys_processing_methodID) ? r_sub01_U_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 14'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_T_addr = ( (|r_sys_processing_methodID) ? r_sub00_T_addr : 14'sh0 ) ;
	assign w_sub00_T_datain = ( (|r_sys_processing_methodID) ? r_sub00_T_datain : 32'h0 ) ;
	assign w_sub00_T_r_w = ( (|r_sys_processing_methodID) ? r_sub00_T_r_w : 1'h0 ) ;
	assign w_sub00_V_addr = ( (|r_sys_processing_methodID) ? r_sub00_V_addr : 14'sh0 ) ;
	assign w_sub00_V_datain = ( (|r_sys_processing_methodID) ? r_sub00_V_datain : 32'h0 ) ;
	assign w_sub00_V_r_w = ( (|r_sys_processing_methodID) ? r_sub00_V_r_w : 1'h0 ) ;
	assign w_sub00_U_addr = ( (|r_sys_processing_methodID) ? r_sub00_U_addr : 14'sh0 ) ;
	assign w_sub00_U_datain = ( (|r_sys_processing_methodID) ? r_sub00_U_datain : 32'h0 ) ;
	assign w_sub00_U_r_w = ( (|r_sys_processing_methodID) ? r_sub00_U_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 14'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub13_T_addr = ( (|r_sys_processing_methodID) ? r_sub13_T_addr : 14'sh0 ) ;
	assign w_sub13_T_datain = ( (|r_sys_processing_methodID) ? r_sub13_T_datain : 32'h0 ) ;
	assign w_sub13_T_r_w = ( (|r_sys_processing_methodID) ? r_sub13_T_r_w : 1'h0 ) ;
	assign w_sub13_V_addr = ( (|r_sys_processing_methodID) ? r_sub13_V_addr : 14'sh0 ) ;
	assign w_sub13_V_datain = ( (|r_sys_processing_methodID) ? r_sub13_V_datain : 32'h0 ) ;
	assign w_sub13_V_r_w = ( (|r_sys_processing_methodID) ? r_sub13_V_r_w : 1'h0 ) ;
	assign w_sub13_U_addr = ( (|r_sys_processing_methodID) ? r_sub13_U_addr : 14'sh0 ) ;
	assign w_sub13_U_datain = ( (|r_sys_processing_methodID) ? r_sub13_U_datain : 32'h0 ) ;
	assign w_sub13_U_r_w = ( (|r_sys_processing_methodID) ? r_sub13_U_r_w : 1'h0 ) ;
	assign w_sub13_result_addr = ( (|r_sys_processing_methodID) ? r_sub13_result_addr : 14'sh0 ) ;
	assign w_sub13_result_datain = ( (|r_sys_processing_methodID) ? r_sub13_result_datain : 32'h0 ) ;
	assign w_sub13_result_r_w = ( (|r_sys_processing_methodID) ? r_sub13_result_r_w : 1'h0 ) ;
	assign w_sub07_T_addr = ( (|r_sys_processing_methodID) ? r_sub07_T_addr : 14'sh0 ) ;
	assign w_sub07_T_datain = ( (|r_sys_processing_methodID) ? r_sub07_T_datain : 32'h0 ) ;
	assign w_sub07_T_r_w = ( (|r_sys_processing_methodID) ? r_sub07_T_r_w : 1'h0 ) ;
	assign w_sub07_V_addr = ( (|r_sys_processing_methodID) ? r_sub07_V_addr : 14'sh0 ) ;
	assign w_sub07_V_datain = ( (|r_sys_processing_methodID) ? r_sub07_V_datain : 32'h0 ) ;
	assign w_sub07_V_r_w = ( (|r_sys_processing_methodID) ? r_sub07_V_r_w : 1'h0 ) ;
	assign w_sub07_U_addr = ( (|r_sys_processing_methodID) ? r_sub07_U_addr : 14'sh0 ) ;
	assign w_sub07_U_datain = ( (|r_sys_processing_methodID) ? r_sub07_U_datain : 32'h0 ) ;
	assign w_sub07_U_r_w = ( (|r_sys_processing_methodID) ? r_sub07_U_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 14'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub16_T_addr = ( (|r_sys_processing_methodID) ? r_sub16_T_addr : 14'sh0 ) ;
	assign w_sub16_T_datain = ( (|r_sys_processing_methodID) ? r_sub16_T_datain : 32'h0 ) ;
	assign w_sub16_T_r_w = ( (|r_sys_processing_methodID) ? r_sub16_T_r_w : 1'h0 ) ;
	assign w_sub16_V_addr = ( (|r_sys_processing_methodID) ? r_sub16_V_addr : 14'sh0 ) ;
	assign w_sub16_V_datain = ( (|r_sys_processing_methodID) ? r_sub16_V_datain : 32'h0 ) ;
	assign w_sub16_V_r_w = ( (|r_sys_processing_methodID) ? r_sub16_V_r_w : 1'h0 ) ;
	assign w_sub16_U_addr = ( (|r_sys_processing_methodID) ? r_sub16_U_addr : 14'sh0 ) ;
	assign w_sub16_U_datain = ( (|r_sys_processing_methodID) ? r_sub16_U_datain : 32'h0 ) ;
	assign w_sub16_U_r_w = ( (|r_sys_processing_methodID) ? r_sub16_U_r_w : 1'h0 ) ;
	assign w_sub16_result_addr = ( (|r_sys_processing_methodID) ? r_sub16_result_addr : 14'sh0 ) ;
	assign w_sub16_result_datain = ( (|r_sys_processing_methodID) ? r_sub16_result_datain : 32'h0 ) ;
	assign w_sub16_result_r_w = ( (|r_sys_processing_methodID) ? r_sub16_result_r_w : 1'h0 ) ;
	assign w_sub06_T_addr = ( (|r_sys_processing_methodID) ? r_sub06_T_addr : 14'sh0 ) ;
	assign w_sub06_T_datain = ( (|r_sys_processing_methodID) ? r_sub06_T_datain : 32'h0 ) ;
	assign w_sub06_T_r_w = ( (|r_sys_processing_methodID) ? r_sub06_T_r_w : 1'h0 ) ;
	assign w_sub06_V_addr = ( (|r_sys_processing_methodID) ? r_sub06_V_addr : 14'sh0 ) ;
	assign w_sub06_V_datain = ( (|r_sys_processing_methodID) ? r_sub06_V_datain : 32'h0 ) ;
	assign w_sub06_V_r_w = ( (|r_sys_processing_methodID) ? r_sub06_V_r_w : 1'h0 ) ;
	assign w_sub06_U_addr = ( (|r_sys_processing_methodID) ? r_sub06_U_addr : 14'sh0 ) ;
	assign w_sub06_U_datain = ( (|r_sys_processing_methodID) ? r_sub06_U_datain : 32'h0 ) ;
	assign w_sub06_U_r_w = ( (|r_sys_processing_methodID) ? r_sub06_U_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 14'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub15_T_addr = ( (|r_sys_processing_methodID) ? r_sub15_T_addr : 14'sh0 ) ;
	assign w_sub15_T_datain = ( (|r_sys_processing_methodID) ? r_sub15_T_datain : 32'h0 ) ;
	assign w_sub15_T_r_w = ( (|r_sys_processing_methodID) ? r_sub15_T_r_w : 1'h0 ) ;
	assign w_sub15_V_addr = ( (|r_sys_processing_methodID) ? r_sub15_V_addr : 14'sh0 ) ;
	assign w_sub15_V_datain = ( (|r_sys_processing_methodID) ? r_sub15_V_datain : 32'h0 ) ;
	assign w_sub15_V_r_w = ( (|r_sys_processing_methodID) ? r_sub15_V_r_w : 1'h0 ) ;
	assign w_sub15_U_addr = ( (|r_sys_processing_methodID) ? r_sub15_U_addr : 14'sh0 ) ;
	assign w_sub15_U_datain = ( (|r_sys_processing_methodID) ? r_sub15_U_datain : 32'h0 ) ;
	assign w_sub15_U_r_w = ( (|r_sys_processing_methodID) ? r_sub15_U_r_w : 1'h0 ) ;
	assign w_sub15_result_addr = ( (|r_sys_processing_methodID) ? r_sub15_result_addr : 14'sh0 ) ;
	assign w_sub15_result_datain = ( (|r_sys_processing_methodID) ? r_sub15_result_datain : 32'h0 ) ;
	assign w_sub15_result_r_w = ( (|r_sys_processing_methodID) ? r_sub15_result_r_w : 1'h0 ) ;
	assign w_sub05_T_addr = ( (|r_sys_processing_methodID) ? r_sub05_T_addr : 14'sh0 ) ;
	assign w_sub05_T_datain = ( (|r_sys_processing_methodID) ? r_sub05_T_datain : 32'h0 ) ;
	assign w_sub05_T_r_w = ( (|r_sys_processing_methodID) ? r_sub05_T_r_w : 1'h0 ) ;
	assign w_sub05_V_addr = ( (|r_sys_processing_methodID) ? r_sub05_V_addr : 14'sh0 ) ;
	assign w_sub05_V_datain = ( (|r_sys_processing_methodID) ? r_sub05_V_datain : 32'h0 ) ;
	assign w_sub05_V_r_w = ( (|r_sys_processing_methodID) ? r_sub05_V_r_w : 1'h0 ) ;
	assign w_sub05_U_addr = ( (|r_sys_processing_methodID) ? r_sub05_U_addr : 14'sh0 ) ;
	assign w_sub05_U_datain = ( (|r_sys_processing_methodID) ? r_sub05_U_datain : 32'h0 ) ;
	assign w_sub05_U_r_w = ( (|r_sys_processing_methodID) ? r_sub05_U_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 14'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub18_T_addr = ( (|r_sys_processing_methodID) ? r_sub18_T_addr : 14'sh0 ) ;
	assign w_sub18_T_datain = ( (|r_sys_processing_methodID) ? r_sub18_T_datain : 32'h0 ) ;
	assign w_sub18_T_r_w = ( (|r_sys_processing_methodID) ? r_sub18_T_r_w : 1'h0 ) ;
	assign w_sub18_V_addr = ( (|r_sys_processing_methodID) ? r_sub18_V_addr : 14'sh0 ) ;
	assign w_sub18_V_datain = ( (|r_sys_processing_methodID) ? r_sub18_V_datain : 32'h0 ) ;
	assign w_sub18_V_r_w = ( (|r_sys_processing_methodID) ? r_sub18_V_r_w : 1'h0 ) ;
	assign w_sub18_U_addr = ( (|r_sys_processing_methodID) ? r_sub18_U_addr : 14'sh0 ) ;
	assign w_sub18_U_datain = ( (|r_sys_processing_methodID) ? r_sub18_U_datain : 32'h0 ) ;
	assign w_sub18_U_r_w = ( (|r_sys_processing_methodID) ? r_sub18_U_r_w : 1'h0 ) ;
	assign w_sub18_result_addr = ( (|r_sys_processing_methodID) ? r_sub18_result_addr : 14'sh0 ) ;
	assign w_sub18_result_datain = ( (|r_sys_processing_methodID) ? r_sub18_result_datain : 32'h0 ) ;
	assign w_sub18_result_r_w = ( (|r_sys_processing_methodID) ? r_sub18_result_r_w : 1'h0 ) ;
	assign w_sub04_T_addr = ( (|r_sys_processing_methodID) ? r_sub04_T_addr : 14'sh0 ) ;
	assign w_sub04_T_datain = ( (|r_sys_processing_methodID) ? r_sub04_T_datain : 32'h0 ) ;
	assign w_sub04_T_r_w = ( (|r_sys_processing_methodID) ? r_sub04_T_r_w : 1'h0 ) ;
	assign w_sub04_V_addr = ( (|r_sys_processing_methodID) ? r_sub04_V_addr : 14'sh0 ) ;
	assign w_sub04_V_datain = ( (|r_sys_processing_methodID) ? r_sub04_V_datain : 32'h0 ) ;
	assign w_sub04_V_r_w = ( (|r_sys_processing_methodID) ? r_sub04_V_r_w : 1'h0 ) ;
	assign w_sub04_U_addr = ( (|r_sys_processing_methodID) ? r_sub04_U_addr : 14'sh0 ) ;
	assign w_sub04_U_datain = ( (|r_sys_processing_methodID) ? r_sub04_U_datain : 32'h0 ) ;
	assign w_sub04_U_r_w = ( (|r_sys_processing_methodID) ? r_sub04_U_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 14'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sub17_T_addr = ( (|r_sys_processing_methodID) ? r_sub17_T_addr : 14'sh0 ) ;
	assign w_sub17_T_datain = ( (|r_sys_processing_methodID) ? r_sub17_T_datain : 32'h0 ) ;
	assign w_sub17_T_r_w = ( (|r_sys_processing_methodID) ? r_sub17_T_r_w : 1'h0 ) ;
	assign w_sub17_V_addr = ( (|r_sys_processing_methodID) ? r_sub17_V_addr : 14'sh0 ) ;
	assign w_sub17_V_datain = ( (|r_sys_processing_methodID) ? r_sub17_V_datain : 32'h0 ) ;
	assign w_sub17_V_r_w = ( (|r_sys_processing_methodID) ? r_sub17_V_r_w : 1'h0 ) ;
	assign w_sub17_U_addr = ( (|r_sys_processing_methodID) ? r_sub17_U_addr : 14'sh0 ) ;
	assign w_sub17_U_datain = ( (|r_sys_processing_methodID) ? r_sub17_U_datain : 32'h0 ) ;
	assign w_sub17_U_r_w = ( (|r_sys_processing_methodID) ? r_sub17_U_r_w : 1'h0 ) ;
	assign w_sub17_result_addr = ( (|r_sys_processing_methodID) ? r_sub17_result_addr : 14'sh0 ) ;
	assign w_sub17_result_datain = ( (|r_sys_processing_methodID) ? r_sub17_result_datain : 32'h0 ) ;
	assign w_sub17_result_r_w = ( (|r_sys_processing_methodID) ? r_sub17_result_r_w : 1'h0 ) ;
	assign w_sub10_T_addr = ( (|r_sys_processing_methodID) ? r_sub10_T_addr : 14'sh0 ) ;
	assign w_sub10_T_datain = ( (|r_sys_processing_methodID) ? r_sub10_T_datain : 32'h0 ) ;
	assign w_sub10_T_r_w = ( (|r_sys_processing_methodID) ? r_sub10_T_r_w : 1'h0 ) ;
	assign w_sub10_V_addr = ( (|r_sys_processing_methodID) ? r_sub10_V_addr : 14'sh0 ) ;
	assign w_sub10_V_datain = ( (|r_sys_processing_methodID) ? r_sub10_V_datain : 32'h0 ) ;
	assign w_sub10_V_r_w = ( (|r_sys_processing_methodID) ? r_sub10_V_r_w : 1'h0 ) ;
	assign w_sub10_U_addr = ( (|r_sys_processing_methodID) ? r_sub10_U_addr : 14'sh0 ) ;
	assign w_sub10_U_datain = ( (|r_sys_processing_methodID) ? r_sub10_U_datain : 32'h0 ) ;
	assign w_sub10_U_r_w = ( (|r_sys_processing_methodID) ? r_sub10_U_r_w : 1'h0 ) ;
	assign w_sub10_result_addr = ( (|r_sys_processing_methodID) ? r_sub10_result_addr : 14'sh0 ) ;
	assign w_sub10_result_datain = ( (|r_sys_processing_methodID) ? r_sub10_result_datain : 32'h0 ) ;
	assign w_sub10_result_r_w = ( (|r_sys_processing_methodID) ? r_sub10_result_r_w : 1'h0 ) ;
	assign w_sub20_T_addr = ( (|r_sys_processing_methodID) ? r_sub20_T_addr : 14'sh0 ) ;
	assign w_sub20_T_datain = ( (|r_sys_processing_methodID) ? r_sub20_T_datain : 32'h0 ) ;
	assign w_sub20_T_r_w = ( (|r_sys_processing_methodID) ? r_sub20_T_r_w : 1'h0 ) ;
	assign w_sub20_V_addr = ( (|r_sys_processing_methodID) ? r_sub20_V_addr : 14'sh0 ) ;
	assign w_sub20_V_datain = ( (|r_sys_processing_methodID) ? r_sub20_V_datain : 32'h0 ) ;
	assign w_sub20_V_r_w = ( (|r_sys_processing_methodID) ? r_sub20_V_r_w : 1'h0 ) ;
	assign w_sub20_U_addr = ( (|r_sys_processing_methodID) ? r_sub20_U_addr : 14'sh0 ) ;
	assign w_sub20_U_datain = ( (|r_sys_processing_methodID) ? r_sub20_U_datain : 32'h0 ) ;
	assign w_sub20_U_r_w = ( (|r_sys_processing_methodID) ? r_sub20_U_r_w : 1'h0 ) ;
	assign w_sub20_result_addr = ( (|r_sys_processing_methodID) ? r_sub20_result_addr : 14'sh0 ) ;
	assign w_sub20_result_datain = ( (|r_sys_processing_methodID) ? r_sub20_result_datain : 32'h0 ) ;
	assign w_sub20_result_r_w = ( (|r_sys_processing_methodID) ? r_sub20_result_r_w : 1'h0 ) ;
	assign w_sub21_T_addr = ( (|r_sys_processing_methodID) ? r_sub21_T_addr : 14'sh0 ) ;
	assign w_sub21_T_datain = ( (|r_sys_processing_methodID) ? r_sub21_T_datain : 32'h0 ) ;
	assign w_sub21_T_r_w = ( (|r_sys_processing_methodID) ? r_sub21_T_r_w : 1'h0 ) ;
	assign w_sub21_V_addr = ( (|r_sys_processing_methodID) ? r_sub21_V_addr : 14'sh0 ) ;
	assign w_sub21_V_datain = ( (|r_sys_processing_methodID) ? r_sub21_V_datain : 32'h0 ) ;
	assign w_sub21_V_r_w = ( (|r_sys_processing_methodID) ? r_sub21_V_r_w : 1'h0 ) ;
	assign w_sub21_U_addr = ( (|r_sys_processing_methodID) ? r_sub21_U_addr : 14'sh0 ) ;
	assign w_sub21_U_datain = ( (|r_sys_processing_methodID) ? r_sub21_U_datain : 32'h0 ) ;
	assign w_sub21_U_r_w = ( (|r_sys_processing_methodID) ? r_sub21_U_r_w : 1'h0 ) ;
	assign w_sub21_result_addr = ( (|r_sys_processing_methodID) ? r_sub21_result_addr : 14'sh0 ) ;
	assign w_sub21_result_datain = ( (|r_sys_processing_methodID) ? r_sub21_result_datain : 32'h0 ) ;
	assign w_sub21_result_r_w = ( (|r_sys_processing_methodID) ? r_sub21_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh00000064;
	assign w_sys_tmp3 = 32'sh00000065;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'h3d23d70a;
	assign w_sys_tmp7 = 32'h3c23d70a;
	assign w_sys_tmp8 = 32'h3bccccce;
	assign w_sys_tmp9 = 32'h3cccccce;
	assign w_sys_tmp10 = 32'h3ea00001;
	assign w_sys_tmp11 = 32'h40a00001;
	assign w_sys_tmp12 = ( !w_sys_tmp13 );
	assign w_sys_tmp13 = (r_run_my_33 < r_run_k_29);
	assign w_sys_tmp14 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp15 = ( !w_sys_tmp16 );
	assign w_sys_tmp16 = (r_run_mx_32 < r_run_j_30);
	assign w_sys_tmp18 = w_ip_MultFloat_product_0;
	assign w_sys_tmp19 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp20 = (r_run_k_29 - w_sys_intOne);
	assign w_sys_tmp22 = (w_sys_tmp23 + r_run_k_29);
	assign w_sys_tmp23 = (r_run_j_30 * w_sys_tmp24);
	assign w_sys_tmp24 = 32'sh00000065;
	assign w_sys_tmp25 = 32'h0;
	assign w_sys_tmp27 = (w_sys_tmp28 + r_run_k_29);
	assign w_sys_tmp28 = (r_run_copy2_j_47 * w_sys_tmp24);
	assign w_sys_tmp32 = (w_sys_tmp33 + r_run_k_29);
	assign w_sys_tmp33 = (r_run_copy1_j_46 * w_sys_tmp24);
	assign w_sys_tmp36 = 32'h42200000;
	assign w_sys_tmp37 = w_sys_tmp18;
	assign w_sys_tmp38 = 32'h3f800000;
	assign w_sys_tmp41 = (w_sys_tmp42 + r_run_k_29);
	assign w_sys_tmp42 = (r_run_copy0_j_45 * w_sys_tmp24);
	assign w_sys_tmp45 = (r_run_copy0_j_45 + w_sys_intOne);
	assign w_sys_tmp46 = (r_run_copy1_j_46 + w_sys_intOne);
	assign w_sys_tmp47 = (r_run_copy2_j_47 + w_sys_intOne);
	assign w_sys_tmp48 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp128 = r_sys_tmp17_float;
	assign w_sys_tmp157 = r_sys_tmp16_float;
	assign w_sys_tmp185 = r_sys_tmp14_float;
	assign w_sys_tmp213 = r_sys_tmp10_float;
	assign w_sys_tmp269 = r_sys_tmp9_float;
	assign w_sys_tmp297 = r_sys_tmp8_float;
	assign w_sys_tmp588 = ( !w_sys_tmp589 );
	assign w_sys_tmp589 = (w_sys_tmp590 < r_run_k_29);
	assign w_sys_tmp590 = 32'sh00000016;
	assign w_sys_tmp593 = (w_sys_tmp594 + r_run_k_29);
	assign w_sys_tmp594 = 32'sh00000065;
	assign w_sys_tmp595 = w_fld_U_2_dataout_1;
	assign w_sys_tmp601 = w_fld_V_3_dataout_1;
	assign w_sys_tmp605 = (w_sys_tmp606 + r_run_k_29);
	assign w_sys_tmp606 = 32'sh000000ca;
	assign w_sys_tmp617 = (w_sys_tmp618 + r_run_k_29);
	assign w_sys_tmp618 = 32'sh0000012f;
	assign w_sys_tmp629 = (w_sys_tmp630 + r_run_k_29);
	assign w_sys_tmp630 = 32'sh00000194;
	assign w_sys_tmp641 = (w_sys_tmp642 + r_run_k_29);
	assign w_sys_tmp642 = 32'sh000001f9;
	assign w_sys_tmp653 = (w_sys_tmp654 + r_run_k_29);
	assign w_sys_tmp654 = 32'sh0000025e;
	assign w_sys_tmp665 = (w_sys_tmp666 + r_run_k_29);
	assign w_sys_tmp666 = 32'sh000002c3;
	assign w_sys_tmp677 = (w_sys_tmp678 + r_run_k_29);
	assign w_sys_tmp678 = 32'sh00000328;
	assign w_sys_tmp689 = (w_sys_tmp690 + r_run_k_29);
	assign w_sys_tmp690 = 32'sh0000038d;
	assign w_sys_tmp701 = (w_sys_tmp702 + r_run_k_29);
	assign w_sys_tmp702 = 32'sh000003f2;
	assign w_sys_tmp713 = (w_sys_tmp714 + r_run_k_29);
	assign w_sys_tmp714 = 32'sh00000457;
	assign w_sys_tmp725 = (w_sys_tmp726 + r_run_k_29);
	assign w_sys_tmp726 = 32'sh000004bc;
	assign w_sys_tmp737 = (w_sys_tmp738 + r_run_k_29);
	assign w_sys_tmp738 = 32'sh00000521;
	assign w_sys_tmp749 = (w_sys_tmp750 + r_run_k_29);
	assign w_sys_tmp750 = 32'sh00000586;
	assign w_sys_tmp761 = (w_sys_tmp762 + r_run_k_29);
	assign w_sys_tmp762 = 32'sh000005eb;
	assign w_sys_tmp773 = (w_sys_tmp774 + r_run_k_29);
	assign w_sys_tmp774 = 32'sh00000650;
	assign w_sys_tmp785 = (w_sys_tmp786 + r_run_k_29);
	assign w_sys_tmp786 = 32'sh000006b5;
	assign w_sys_tmp797 = (w_sys_tmp798 + r_run_k_29);
	assign w_sys_tmp798 = 32'sh0000071a;
	assign w_sys_tmp809 = (w_sys_tmp810 + r_run_k_29);
	assign w_sys_tmp810 = 32'sh0000077f;
	assign w_sys_tmp821 = (w_sys_tmp822 + r_run_k_29);
	assign w_sys_tmp822 = 32'sh000007e4;
	assign w_sys_tmp833 = (w_sys_tmp834 + r_run_k_29);
	assign w_sys_tmp834 = 32'sh00000849;
	assign w_sys_tmp845 = (w_sys_tmp846 + r_run_k_29);
	assign w_sys_tmp846 = 32'sh000008ae;
	assign w_sys_tmp881 = (w_sys_tmp882 + r_run_k_29);
	assign w_sys_tmp882 = 32'sh00000913;
	assign w_sys_tmp893 = (w_sys_tmp894 + r_run_k_29);
	assign w_sys_tmp894 = 32'sh00000978;
	assign w_sys_tmp905 = (w_sys_tmp906 + r_run_k_29);
	assign w_sys_tmp906 = 32'sh000009dd;
	assign w_sys_tmp917 = (w_sys_tmp918 + r_run_k_29);
	assign w_sys_tmp918 = 32'sh00000a42;
	assign w_sys_tmp929 = (w_sys_tmp930 + r_run_k_29);
	assign w_sys_tmp930 = 32'sh00000aa7;
	assign w_sys_tmp941 = (w_sys_tmp942 + r_run_k_29);
	assign w_sys_tmp942 = 32'sh00000b0c;
	assign w_sys_tmp953 = (w_sys_tmp954 + r_run_k_29);
	assign w_sys_tmp954 = 32'sh00000b71;
	assign w_sys_tmp965 = (w_sys_tmp966 + r_run_k_29);
	assign w_sys_tmp966 = 32'sh00000bd6;
	assign w_sys_tmp977 = (w_sys_tmp978 + r_run_k_29);
	assign w_sys_tmp978 = 32'sh00000c3b;
	assign w_sys_tmp989 = (w_sys_tmp990 + r_run_k_29);
	assign w_sys_tmp990 = 32'sh00000ca0;
	assign w_sys_tmp1001 = (w_sys_tmp1002 + r_run_k_29);
	assign w_sys_tmp1002 = 32'sh00000d05;
	assign w_sys_tmp1013 = (w_sys_tmp1014 + r_run_k_29);
	assign w_sys_tmp1014 = 32'sh00000d6a;
	assign w_sys_tmp1025 = (w_sys_tmp1026 + r_run_k_29);
	assign w_sys_tmp1026 = 32'sh00000dcf;
	assign w_sys_tmp1037 = (w_sys_tmp1038 + r_run_k_29);
	assign w_sys_tmp1038 = 32'sh00000e34;
	assign w_sys_tmp1049 = (w_sys_tmp1050 + r_run_k_29);
	assign w_sys_tmp1050 = 32'sh00000e99;
	assign w_sys_tmp1061 = (w_sys_tmp1062 + r_run_k_29);
	assign w_sys_tmp1062 = 32'sh00000efe;
	assign w_sys_tmp1073 = (w_sys_tmp1074 + r_run_k_29);
	assign w_sys_tmp1074 = 32'sh00000f63;
	assign w_sys_tmp1085 = (w_sys_tmp1086 + r_run_k_29);
	assign w_sys_tmp1086 = 32'sh00000fc8;
	assign w_sys_tmp1097 = (w_sys_tmp1098 + r_run_k_29);
	assign w_sys_tmp1098 = 32'sh0000102d;
	assign w_sys_tmp1109 = (w_sys_tmp1110 + r_run_k_29);
	assign w_sys_tmp1110 = 32'sh00001092;
	assign w_sys_tmp1145 = (w_sys_tmp1146 + r_run_k_29);
	assign w_sys_tmp1146 = 32'sh000010f7;
	assign w_sys_tmp1157 = (w_sys_tmp1158 + r_run_k_29);
	assign w_sys_tmp1158 = 32'sh0000115c;
	assign w_sys_tmp1169 = (w_sys_tmp1170 + r_run_k_29);
	assign w_sys_tmp1170 = 32'sh000011c1;
	assign w_sys_tmp1181 = (w_sys_tmp1182 + r_run_k_29);
	assign w_sys_tmp1182 = 32'sh00001226;
	assign w_sys_tmp1193 = (w_sys_tmp1194 + r_run_k_29);
	assign w_sys_tmp1194 = 32'sh0000128b;
	assign w_sys_tmp1205 = (w_sys_tmp1206 + r_run_k_29);
	assign w_sys_tmp1206 = 32'sh00019670;
	assign w_sys_tmp1217 = (w_sys_tmp1218 + r_run_k_29);
	assign w_sys_tmp1218 = 32'sh00001355;
	assign w_sys_tmp1229 = (w_sys_tmp1230 + r_run_k_29);
	assign w_sys_tmp1230 = 32'sh000013ba;
	assign w_sys_tmp1241 = (w_sys_tmp1242 + r_run_k_29);
	assign w_sys_tmp1242 = 32'sh0000141f;
	assign w_sys_tmp1253 = (w_sys_tmp1254 + r_run_k_29);
	assign w_sys_tmp1254 = 32'sh00001484;
	assign w_sys_tmp1265 = (w_sys_tmp1266 + r_run_k_29);
	assign w_sys_tmp1266 = 32'sh000014e9;
	assign w_sys_tmp1277 = (w_sys_tmp1278 + r_run_k_29);
	assign w_sys_tmp1278 = 32'sh0000154e;
	assign w_sys_tmp1289 = (w_sys_tmp1290 + r_run_k_29);
	assign w_sys_tmp1290 = 32'sh000015b3;
	assign w_sys_tmp1301 = (w_sys_tmp1302 + r_run_k_29);
	assign w_sys_tmp1302 = 32'sh00001618;
	assign w_sys_tmp1313 = (w_sys_tmp1314 + r_run_k_29);
	assign w_sys_tmp1314 = 32'sh0000167d;
	assign w_sys_tmp1325 = (w_sys_tmp1326 + r_run_k_29);
	assign w_sys_tmp1326 = 32'sh000016e2;
	assign w_sys_tmp1337 = (w_sys_tmp1338 + r_run_k_29);
	assign w_sys_tmp1338 = 32'sh00001747;
	assign w_sys_tmp1349 = (w_sys_tmp1350 + r_run_k_29);
	assign w_sys_tmp1350 = 32'sh000017ac;
	assign w_sys_tmp1361 = (w_sys_tmp1362 + r_run_k_29);
	assign w_sys_tmp1362 = 32'sh00001811;
	assign w_sys_tmp1385 = (w_sys_tmp1386 + r_run_k_29);
	assign w_sys_tmp1386 = 32'sh00001876;
	assign w_sys_tmp1397 = (w_sys_tmp1398 + r_run_k_29);
	assign w_sys_tmp1398 = 32'sh000018db;
	assign w_sys_tmp1409 = (w_sys_tmp1410 + r_run_k_29);
	assign w_sys_tmp1410 = 32'sh00001940;
	assign w_sys_tmp1421 = (w_sys_tmp1422 + r_run_k_29);
	assign w_sys_tmp1422 = 32'sh000019a5;
	assign w_sys_tmp1433 = (w_sys_tmp1434 + r_run_k_29);
	assign w_sys_tmp1434 = 32'sh00001a0a;
	assign w_sys_tmp1445 = (w_sys_tmp1446 + r_run_k_29);
	assign w_sys_tmp1446 = 32'sh00001a6f;
	assign w_sys_tmp1457 = (w_sys_tmp1458 + r_run_k_29);
	assign w_sys_tmp1458 = 32'sh00001ad4;
	assign w_sys_tmp1469 = (w_sys_tmp1470 + r_run_k_29);
	assign w_sys_tmp1470 = 32'sh00001b39;
	assign w_sys_tmp1481 = (w_sys_tmp1482 + r_run_k_29);
	assign w_sys_tmp1482 = 32'sh00001b9e;
	assign w_sys_tmp1493 = (w_sys_tmp1494 + r_run_k_29);
	assign w_sys_tmp1494 = 32'sh00001c03;
	assign w_sys_tmp1505 = (w_sys_tmp1506 + r_run_k_29);
	assign w_sys_tmp1506 = 32'sh00001c68;
	assign w_sys_tmp1517 = (w_sys_tmp1518 + r_run_k_29);
	assign w_sys_tmp1518 = 32'sh00001ccd;
	assign w_sys_tmp1529 = (w_sys_tmp1530 + r_run_k_29);
	assign w_sys_tmp1530 = 32'sh00001d32;
	assign w_sys_tmp1541 = (w_sys_tmp1542 + r_run_k_29);
	assign w_sys_tmp1542 = 32'sh00001d97;
	assign w_sys_tmp1553 = (w_sys_tmp1554 + r_run_k_29);
	assign w_sys_tmp1554 = 32'sh00001dfc;
	assign w_sys_tmp1565 = (w_sys_tmp1566 + r_run_k_29);
	assign w_sys_tmp1566 = 32'sh00001e61;
	assign w_sys_tmp1577 = (w_sys_tmp1578 + r_run_k_29);
	assign w_sys_tmp1578 = 32'sh00001ec6;
	assign w_sys_tmp1589 = (w_sys_tmp1590 + r_run_k_29);
	assign w_sys_tmp1590 = 32'sh00001f2b;
	assign w_sys_tmp1601 = (w_sys_tmp1602 + r_run_k_29);
	assign w_sys_tmp1602 = 32'sh00001f90;
	assign w_sys_tmp1613 = (w_sys_tmp1614 + r_run_k_29);
	assign w_sys_tmp1614 = 32'sh00001ff5;
	assign w_sys_tmp1625 = (w_sys_tmp1626 + r_run_k_29);
	assign w_sys_tmp1626 = 32'sh0000205a;
	assign w_sys_tmp1661 = (w_sys_tmp1662 + r_run_k_29);
	assign w_sys_tmp1662 = 32'sh000020bf;
	assign w_sys_tmp1673 = (w_sys_tmp1674 + r_run_k_29);
	assign w_sys_tmp1674 = 32'sh000c5da4;
	assign w_sys_tmp1685 = (w_sys_tmp1686 + r_run_k_29);
	assign w_sys_tmp1686 = 32'sh00002189;
	assign w_sys_tmp1697 = (w_sys_tmp1698 + r_run_k_29);
	assign w_sys_tmp1698 = 32'sh000021ee;
	assign w_sys_tmp1709 = (w_sys_tmp1710 + r_run_k_29);
	assign w_sys_tmp1710 = 32'sh00002253;
	assign w_sys_tmp1721 = (w_sys_tmp1722 + r_run_k_29);
	assign w_sys_tmp1722 = 32'sh000022b8;
	assign w_sys_tmp1733 = (w_sys_tmp1734 + r_run_k_29);
	assign w_sys_tmp1734 = 32'sh0000231d;
	assign w_sys_tmp1745 = (w_sys_tmp1746 + r_run_k_29);
	assign w_sys_tmp1746 = 32'sh00002382;
	assign w_sys_tmp1757 = (w_sys_tmp1758 + r_run_k_29);
	assign w_sys_tmp1758 = 32'sh000023e7;
	assign w_sys_tmp1769 = (w_sys_tmp1770 + r_run_k_29);
	assign w_sys_tmp1770 = 32'sh0000244c;
	assign w_sys_tmp1781 = (w_sys_tmp1782 + r_run_k_29);
	assign w_sys_tmp1782 = 32'sh000024b1;
	assign w_sys_tmp1793 = (w_sys_tmp1794 + r_run_k_29);
	assign w_sys_tmp1794 = 32'sh00002516;
	assign w_sys_tmp1805 = (w_sys_tmp1806 + r_run_k_29);
	assign w_sys_tmp1806 = 32'sh0000257b;
	assign w_sys_tmp1817 = (w_sys_tmp1818 + r_run_k_29);
	assign w_sys_tmp1818 = 32'sh000025e0;
	assign w_sys_tmp1829 = (w_sys_tmp1830 + r_run_k_29);
	assign w_sys_tmp1830 = 32'sh00002645;
	assign w_sys_tmp1841 = (w_sys_tmp1842 + r_run_k_29);
	assign w_sys_tmp1842 = 32'sh000026aa;
	assign w_sys_tmp1853 = (w_sys_tmp1854 + r_run_k_29);
	assign w_sys_tmp1854 = 32'sh0000270f;
	assign w_sys_tmp1865 = (w_sys_tmp1866 + r_run_k_29);
	assign w_sys_tmp1866 = 32'sh00002774;
	assign w_sys_tmp1877 = (w_sys_tmp1878 + r_run_k_29);
	assign w_sys_tmp1878 = 32'sh000027d9;
	assign w_sys_tmp1889 = (w_sys_tmp1890 + r_run_k_29);
	assign w_sys_tmp1890 = 32'sh00000079;
	assign w_sys_tmp1901 = (w_sys_tmp1902 + r_run_k_29);
	assign w_sys_tmp1902 = 32'sh000000de;
	assign w_sys_tmp1913 = (w_sys_tmp1914 + r_run_k_29);
	assign w_sys_tmp1914 = 32'sh00000143;
	assign w_sys_tmp1925 = (w_sys_tmp1926 + r_run_k_29);
	assign w_sys_tmp1926 = 32'sh000001a8;
	assign w_sys_tmp1937 = (w_sys_tmp1938 + r_run_k_29);
	assign w_sys_tmp1938 = 32'sh0000020d;
	assign w_sys_tmp1949 = (w_sys_tmp1950 + r_run_k_29);
	assign w_sys_tmp1950 = 32'sh00000272;
	assign w_sys_tmp1961 = (w_sys_tmp1962 + r_run_k_29);
	assign w_sys_tmp1962 = 32'sh000002d7;
	assign w_sys_tmp1973 = (w_sys_tmp1974 + r_run_k_29);
	assign w_sys_tmp1974 = 32'sh0000033c;
	assign w_sys_tmp1985 = (w_sys_tmp1986 + r_run_k_29);
	assign w_sys_tmp1986 = 32'sh000003a1;
	assign w_sys_tmp1997 = (w_sys_tmp1998 + r_run_k_29);
	assign w_sys_tmp1998 = 32'sh00000406;
	assign w_sys_tmp2009 = (w_sys_tmp2010 + r_run_k_29);
	assign w_sys_tmp2010 = 32'sh0000046b;
	assign w_sys_tmp2021 = (w_sys_tmp2022 + r_run_k_29);
	assign w_sys_tmp2022 = 32'sh000004d0;
	assign w_sys_tmp2033 = (w_sys_tmp2034 + r_run_k_29);
	assign w_sys_tmp2034 = 32'sh00000535;
	assign w_sys_tmp2045 = (w_sys_tmp2046 + r_run_k_29);
	assign w_sys_tmp2046 = 32'sh0000059a;
	assign w_sys_tmp2057 = (w_sys_tmp2058 + r_run_k_29);
	assign w_sys_tmp2058 = 32'sh000005ff;
	assign w_sys_tmp2069 = (w_sys_tmp2070 + r_run_k_29);
	assign w_sys_tmp2070 = 32'sh00000664;
	assign w_sys_tmp2081 = (w_sys_tmp2082 + r_run_k_29);
	assign w_sys_tmp2082 = 32'sh000006c9;
	assign w_sys_tmp2093 = (w_sys_tmp2094 + r_run_k_29);
	assign w_sys_tmp2094 = 32'sh0000072e;
	assign w_sys_tmp2105 = (w_sys_tmp2106 + r_run_k_29);
	assign w_sys_tmp2106 = 32'sh00000793;
	assign w_sys_tmp2117 = (w_sys_tmp2118 + r_run_k_29);
	assign w_sys_tmp2118 = 32'sh000007f8;
	assign w_sys_tmp2129 = (w_sys_tmp2130 + r_run_k_29);
	assign w_sys_tmp2130 = 32'sh0000085d;
	assign w_sys_tmp2153 = (w_sys_tmp2154 + r_run_k_29);
	assign w_sys_tmp2154 = 32'sh000008c2;
	assign w_sys_tmp2165 = (w_sys_tmp2166 + r_run_k_29);
	assign w_sys_tmp2166 = 32'sh00000927;
	assign w_sys_tmp2177 = (w_sys_tmp2178 + r_run_k_29);
	assign w_sys_tmp2178 = 32'sh0000098c;
	assign w_sys_tmp2189 = (w_sys_tmp2190 + r_run_k_29);
	assign w_sys_tmp2190 = 32'sh000009f1;
	assign w_sys_tmp2201 = (w_sys_tmp2202 + r_run_k_29);
	assign w_sys_tmp2202 = 32'sh00000a56;
	assign w_sys_tmp2213 = (w_sys_tmp2214 + r_run_k_29);
	assign w_sys_tmp2214 = 32'sh00000abb;
	assign w_sys_tmp2225 = (w_sys_tmp2226 + r_run_k_29);
	assign w_sys_tmp2226 = 32'sh00000b20;
	assign w_sys_tmp2237 = (w_sys_tmp2238 + r_run_k_29);
	assign w_sys_tmp2238 = 32'sh00000b85;
	assign w_sys_tmp2249 = (w_sys_tmp2250 + r_run_k_29);
	assign w_sys_tmp2250 = 32'sh00000bea;
	assign w_sys_tmp2261 = (w_sys_tmp2262 + r_run_k_29);
	assign w_sys_tmp2262 = 32'sh00000c4f;
	assign w_sys_tmp2273 = (w_sys_tmp2274 + r_run_k_29);
	assign w_sys_tmp2274 = 32'sh00000cb4;
	assign w_sys_tmp2285 = (w_sys_tmp2286 + r_run_k_29);
	assign w_sys_tmp2286 = 32'sh00000d19;
	assign w_sys_tmp2297 = (w_sys_tmp2298 + r_run_k_29);
	assign w_sys_tmp2298 = 32'sh00000d7e;
	assign w_sys_tmp2309 = (w_sys_tmp2310 + r_run_k_29);
	assign w_sys_tmp2310 = 32'sh00000de3;
	assign w_sys_tmp2321 = (w_sys_tmp2322 + r_run_k_29);
	assign w_sys_tmp2322 = 32'sh00000e48;
	assign w_sys_tmp2333 = (w_sys_tmp2334 + r_run_k_29);
	assign w_sys_tmp2334 = 32'sh00000ead;
	assign w_sys_tmp2345 = (w_sys_tmp2346 + r_run_k_29);
	assign w_sys_tmp2346 = 32'sh00000f12;
	assign w_sys_tmp2357 = (w_sys_tmp2358 + r_run_k_29);
	assign w_sys_tmp2358 = 32'sh00000f77;
	assign w_sys_tmp2369 = (w_sys_tmp2370 + r_run_k_29);
	assign w_sys_tmp2370 = 32'sh00000fdc;
	assign w_sys_tmp2381 = (w_sys_tmp2382 + r_run_k_29);
	assign w_sys_tmp2382 = 32'sh00001041;
	assign w_sys_tmp2393 = (w_sys_tmp2394 + r_run_k_29);
	assign w_sys_tmp2394 = 32'sh000010a6;
	assign w_sys_tmp2429 = (w_sys_tmp2430 + r_run_k_29);
	assign w_sys_tmp2430 = 32'sh0000110b;
	assign w_sys_tmp2441 = (w_sys_tmp2442 + r_run_k_29);
	assign w_sys_tmp2442 = 32'sh00001170;
	assign w_sys_tmp2453 = (w_sys_tmp2454 + r_run_k_29);
	assign w_sys_tmp2454 = 32'sh000011d5;
	assign w_sys_tmp2465 = (w_sys_tmp2466 + r_run_k_29);
	assign w_sys_tmp2466 = 32'sh0000123a;
	assign w_sys_tmp2477 = (w_sys_tmp2478 + r_run_k_29);
	assign w_sys_tmp2478 = 32'sh0000129f;
	assign w_sys_tmp2489 = (w_sys_tmp2490 + r_run_k_29);
	assign w_sys_tmp2490 = 32'sh00019684;
	assign w_sys_tmp2501 = (w_sys_tmp2502 + r_run_k_29);
	assign w_sys_tmp2502 = 32'sh00001369;
	assign w_sys_tmp2513 = (w_sys_tmp2514 + r_run_k_29);
	assign w_sys_tmp2514 = 32'sh000013ce;
	assign w_sys_tmp2525 = (w_sys_tmp2526 + r_run_k_29);
	assign w_sys_tmp2526 = 32'sh00001433;
	assign w_sys_tmp2537 = (w_sys_tmp2538 + r_run_k_29);
	assign w_sys_tmp2538 = 32'sh00001498;
	assign w_sys_tmp2549 = (w_sys_tmp2550 + r_run_k_29);
	assign w_sys_tmp2550 = 32'sh000014fd;
	assign w_sys_tmp2561 = (w_sys_tmp2562 + r_run_k_29);
	assign w_sys_tmp2562 = 32'sh00001562;
	assign w_sys_tmp2573 = (w_sys_tmp2574 + r_run_k_29);
	assign w_sys_tmp2574 = 32'sh000015c7;
	assign w_sys_tmp2585 = (w_sys_tmp2586 + r_run_k_29);
	assign w_sys_tmp2586 = 32'sh0000162c;
	assign w_sys_tmp2597 = (w_sys_tmp2598 + r_run_k_29);
	assign w_sys_tmp2598 = 32'sh00001691;
	assign w_sys_tmp2609 = (w_sys_tmp2610 + r_run_k_29);
	assign w_sys_tmp2610 = 32'sh000016f6;
	assign w_sys_tmp2621 = (w_sys_tmp2622 + r_run_k_29);
	assign w_sys_tmp2622 = 32'sh0000175b;
	assign w_sys_tmp2633 = (w_sys_tmp2634 + r_run_k_29);
	assign w_sys_tmp2634 = 32'sh000017c0;
	assign w_sys_tmp2645 = (w_sys_tmp2646 + r_run_k_29);
	assign w_sys_tmp2646 = 32'sh00001825;
	assign w_sys_tmp2657 = (w_sys_tmp2658 + r_run_k_29);
	assign w_sys_tmp2658 = 32'sh0000188a;
	assign w_sys_tmp2681 = (w_sys_tmp2682 + r_run_k_29);
	assign w_sys_tmp2682 = 32'sh000018ef;
	assign w_sys_tmp2693 = (w_sys_tmp2694 + r_run_k_29);
	assign w_sys_tmp2694 = 32'sh00001954;
	assign w_sys_tmp2705 = (w_sys_tmp2706 + r_run_k_29);
	assign w_sys_tmp2706 = 32'sh000019b9;
	assign w_sys_tmp2717 = (w_sys_tmp2718 + r_run_k_29);
	assign w_sys_tmp2718 = 32'sh00001a1e;
	assign w_sys_tmp2729 = (w_sys_tmp2730 + r_run_k_29);
	assign w_sys_tmp2730 = 32'sh00001a83;
	assign w_sys_tmp2741 = (w_sys_tmp2742 + r_run_k_29);
	assign w_sys_tmp2742 = 32'sh00001ae8;
	assign w_sys_tmp2753 = (w_sys_tmp2754 + r_run_k_29);
	assign w_sys_tmp2754 = 32'sh00001b4d;
	assign w_sys_tmp2765 = (w_sys_tmp2766 + r_run_k_29);
	assign w_sys_tmp2766 = 32'sh00001bb2;
	assign w_sys_tmp2777 = (w_sys_tmp2778 + r_run_k_29);
	assign w_sys_tmp2778 = 32'sh00001c17;
	assign w_sys_tmp2789 = (w_sys_tmp2790 + r_run_k_29);
	assign w_sys_tmp2790 = 32'sh00001c7c;
	assign w_sys_tmp2801 = (w_sys_tmp2802 + r_run_k_29);
	assign w_sys_tmp2802 = 32'sh00001ce1;
	assign w_sys_tmp2813 = (w_sys_tmp2814 + r_run_k_29);
	assign w_sys_tmp2814 = 32'sh00001d46;
	assign w_sys_tmp2825 = (w_sys_tmp2826 + r_run_k_29);
	assign w_sys_tmp2826 = 32'sh00001dab;
	assign w_sys_tmp2837 = (w_sys_tmp2838 + r_run_k_29);
	assign w_sys_tmp2838 = 32'sh00001e10;
	assign w_sys_tmp2849 = (w_sys_tmp2850 + r_run_k_29);
	assign w_sys_tmp2850 = 32'sh00001e75;
	assign w_sys_tmp2861 = (w_sys_tmp2862 + r_run_k_29);
	assign w_sys_tmp2862 = 32'sh00001eda;
	assign w_sys_tmp2873 = (w_sys_tmp2874 + r_run_k_29);
	assign w_sys_tmp2874 = 32'sh00001f3f;
	assign w_sys_tmp2885 = (w_sys_tmp2886 + r_run_k_29);
	assign w_sys_tmp2886 = 32'sh00001fa4;
	assign w_sys_tmp2897 = (w_sys_tmp2898 + r_run_k_29);
	assign w_sys_tmp2898 = 32'sh00002009;
	assign w_sys_tmp2909 = (w_sys_tmp2910 + r_run_k_29);
	assign w_sys_tmp2910 = 32'sh0000206e;
	assign w_sys_tmp2945 = (w_sys_tmp2946 + r_run_k_29);
	assign w_sys_tmp2946 = 32'sh000020d3;
	assign w_sys_tmp2957 = (w_sys_tmp2958 + r_run_k_29);
	assign w_sys_tmp2958 = 32'sh000c5db8;
	assign w_sys_tmp2969 = (w_sys_tmp2970 + r_run_k_29);
	assign w_sys_tmp2970 = 32'sh0000219d;
	assign w_sys_tmp2981 = (w_sys_tmp2982 + r_run_k_29);
	assign w_sys_tmp2982 = 32'sh00002202;
	assign w_sys_tmp2993 = (w_sys_tmp2994 + r_run_k_29);
	assign w_sys_tmp2994 = 32'sh00002267;
	assign w_sys_tmp3005 = (w_sys_tmp3006 + r_run_k_29);
	assign w_sys_tmp3006 = 32'sh000022cc;
	assign w_sys_tmp3017 = (w_sys_tmp3018 + r_run_k_29);
	assign w_sys_tmp3018 = 32'sh00002331;
	assign w_sys_tmp3029 = (w_sys_tmp3030 + r_run_k_29);
	assign w_sys_tmp3030 = 32'sh00002396;
	assign w_sys_tmp3041 = (w_sys_tmp3042 + r_run_k_29);
	assign w_sys_tmp3042 = 32'sh000023fb;
	assign w_sys_tmp3053 = (w_sys_tmp3054 + r_run_k_29);
	assign w_sys_tmp3054 = 32'sh00002460;
	assign w_sys_tmp3065 = (w_sys_tmp3066 + r_run_k_29);
	assign w_sys_tmp3066 = 32'sh000024c5;
	assign w_sys_tmp3077 = (w_sys_tmp3078 + r_run_k_29);
	assign w_sys_tmp3078 = 32'sh0000252a;
	assign w_sys_tmp3089 = (w_sys_tmp3090 + r_run_k_29);
	assign w_sys_tmp3090 = 32'sh0000258f;
	assign w_sys_tmp3101 = (w_sys_tmp3102 + r_run_k_29);
	assign w_sys_tmp3102 = 32'sh000025f4;
	assign w_sys_tmp3113 = (w_sys_tmp3114 + r_run_k_29);
	assign w_sys_tmp3114 = 32'sh00002659;
	assign w_sys_tmp3125 = (w_sys_tmp3126 + r_run_k_29);
	assign w_sys_tmp3126 = 32'sh000026be;
	assign w_sys_tmp3137 = (w_sys_tmp3138 + r_run_k_29);
	assign w_sys_tmp3138 = 32'sh00002723;
	assign w_sys_tmp3149 = (w_sys_tmp3150 + r_run_k_29);
	assign w_sys_tmp3150 = 32'sh00002788;
	assign w_sys_tmp3161 = (w_sys_tmp3162 + r_run_k_29);
	assign w_sys_tmp3162 = 32'sh000027ed;
	assign w_sys_tmp3173 = (w_sys_tmp3174 + r_run_k_29);
	assign w_sys_tmp3174 = 32'sh0000008d;
	assign w_sys_tmp3185 = (w_sys_tmp3186 + r_run_k_29);
	assign w_sys_tmp3186 = 32'sh000000f2;
	assign w_sys_tmp3197 = (w_sys_tmp3198 + r_run_k_29);
	assign w_sys_tmp3198 = 32'sh00000157;
	assign w_sys_tmp3209 = (w_sys_tmp3210 + r_run_k_29);
	assign w_sys_tmp3210 = 32'sh000001bc;
	assign w_sys_tmp3221 = (w_sys_tmp3222 + r_run_k_29);
	assign w_sys_tmp3222 = 32'sh00000221;
	assign w_sys_tmp3233 = (w_sys_tmp3234 + r_run_k_29);
	assign w_sys_tmp3234 = 32'sh00000286;
	assign w_sys_tmp3245 = (w_sys_tmp3246 + r_run_k_29);
	assign w_sys_tmp3246 = 32'sh000002eb;
	assign w_sys_tmp3257 = (w_sys_tmp3258 + r_run_k_29);
	assign w_sys_tmp3258 = 32'sh00000350;
	assign w_sys_tmp3269 = (w_sys_tmp3270 + r_run_k_29);
	assign w_sys_tmp3270 = 32'sh000003b5;
	assign w_sys_tmp3281 = (w_sys_tmp3282 + r_run_k_29);
	assign w_sys_tmp3282 = 32'sh0000041a;
	assign w_sys_tmp3293 = (w_sys_tmp3294 + r_run_k_29);
	assign w_sys_tmp3294 = 32'sh0000047f;
	assign w_sys_tmp3305 = (w_sys_tmp3306 + r_run_k_29);
	assign w_sys_tmp3306 = 32'sh000004e4;
	assign w_sys_tmp3317 = (w_sys_tmp3318 + r_run_k_29);
	assign w_sys_tmp3318 = 32'sh00000549;
	assign w_sys_tmp3329 = (w_sys_tmp3330 + r_run_k_29);
	assign w_sys_tmp3330 = 32'sh000005ae;
	assign w_sys_tmp3341 = (w_sys_tmp3342 + r_run_k_29);
	assign w_sys_tmp3342 = 32'sh00000613;
	assign w_sys_tmp3353 = (w_sys_tmp3354 + r_run_k_29);
	assign w_sys_tmp3354 = 32'sh00000678;
	assign w_sys_tmp3365 = (w_sys_tmp3366 + r_run_k_29);
	assign w_sys_tmp3366 = 32'sh000006dd;
	assign w_sys_tmp3377 = (w_sys_tmp3378 + r_run_k_29);
	assign w_sys_tmp3378 = 32'sh00000742;
	assign w_sys_tmp3389 = (w_sys_tmp3390 + r_run_k_29);
	assign w_sys_tmp3390 = 32'sh000007a7;
	assign w_sys_tmp3401 = (w_sys_tmp3402 + r_run_k_29);
	assign w_sys_tmp3402 = 32'sh0000080c;
	assign w_sys_tmp3413 = (w_sys_tmp3414 + r_run_k_29);
	assign w_sys_tmp3414 = 32'sh00000871;
	assign w_sys_tmp3437 = (w_sys_tmp3438 + r_run_k_29);
	assign w_sys_tmp3438 = 32'sh000008d6;
	assign w_sys_tmp3449 = (w_sys_tmp3450 + r_run_k_29);
	assign w_sys_tmp3450 = 32'sh0000093b;
	assign w_sys_tmp3461 = (w_sys_tmp3462 + r_run_k_29);
	assign w_sys_tmp3462 = 32'sh000009a0;
	assign w_sys_tmp3473 = (w_sys_tmp3474 + r_run_k_29);
	assign w_sys_tmp3474 = 32'sh00000a05;
	assign w_sys_tmp3485 = (w_sys_tmp3486 + r_run_k_29);
	assign w_sys_tmp3486 = 32'sh00000a6a;
	assign w_sys_tmp3497 = (w_sys_tmp3498 + r_run_k_29);
	assign w_sys_tmp3498 = 32'sh00000acf;
	assign w_sys_tmp3509 = (w_sys_tmp3510 + r_run_k_29);
	assign w_sys_tmp3510 = 32'sh00000b34;
	assign w_sys_tmp3521 = (w_sys_tmp3522 + r_run_k_29);
	assign w_sys_tmp3522 = 32'sh00000b99;
	assign w_sys_tmp3533 = (w_sys_tmp3534 + r_run_k_29);
	assign w_sys_tmp3534 = 32'sh00000bfe;
	assign w_sys_tmp3545 = (w_sys_tmp3546 + r_run_k_29);
	assign w_sys_tmp3546 = 32'sh00000c63;
	assign w_sys_tmp3557 = (w_sys_tmp3558 + r_run_k_29);
	assign w_sys_tmp3558 = 32'sh00000cc8;
	assign w_sys_tmp3569 = (w_sys_tmp3570 + r_run_k_29);
	assign w_sys_tmp3570 = 32'sh00000d2d;
	assign w_sys_tmp3581 = (w_sys_tmp3582 + r_run_k_29);
	assign w_sys_tmp3582 = 32'sh00000d92;
	assign w_sys_tmp3593 = (w_sys_tmp3594 + r_run_k_29);
	assign w_sys_tmp3594 = 32'sh00000df7;
	assign w_sys_tmp3605 = (w_sys_tmp3606 + r_run_k_29);
	assign w_sys_tmp3606 = 32'sh00000e5c;
	assign w_sys_tmp3617 = (w_sys_tmp3618 + r_run_k_29);
	assign w_sys_tmp3618 = 32'sh00000ec1;
	assign w_sys_tmp3629 = (w_sys_tmp3630 + r_run_k_29);
	assign w_sys_tmp3630 = 32'sh00000f26;
	assign w_sys_tmp3641 = (w_sys_tmp3642 + r_run_k_29);
	assign w_sys_tmp3642 = 32'sh00000f8b;
	assign w_sys_tmp3653 = (w_sys_tmp3654 + r_run_k_29);
	assign w_sys_tmp3654 = 32'sh00000ff0;
	assign w_sys_tmp3665 = (w_sys_tmp3666 + r_run_k_29);
	assign w_sys_tmp3666 = 32'sh00001055;
	assign w_sys_tmp3677 = (w_sys_tmp3678 + r_run_k_29);
	assign w_sys_tmp3678 = 32'sh000010ba;
	assign w_sys_tmp3713 = (w_sys_tmp3714 + r_run_k_29);
	assign w_sys_tmp3714 = 32'sh0000111f;
	assign w_sys_tmp3725 = (w_sys_tmp3726 + r_run_k_29);
	assign w_sys_tmp3726 = 32'sh00001184;
	assign w_sys_tmp3737 = (w_sys_tmp3738 + r_run_k_29);
	assign w_sys_tmp3738 = 32'sh000011e9;
	assign w_sys_tmp3749 = (w_sys_tmp3750 + r_run_k_29);
	assign w_sys_tmp3750 = 32'sh0000124e;
	assign w_sys_tmp3761 = (w_sys_tmp3762 + r_run_k_29);
	assign w_sys_tmp3762 = 32'sh000012b3;
	assign w_sys_tmp3773 = (w_sys_tmp3774 + r_run_k_29);
	assign w_sys_tmp3774 = 32'sh00019698;
	assign w_sys_tmp3785 = (w_sys_tmp3786 + r_run_k_29);
	assign w_sys_tmp3786 = 32'sh0000137d;
	assign w_sys_tmp3797 = (w_sys_tmp3798 + r_run_k_29);
	assign w_sys_tmp3798 = 32'sh000013e2;
	assign w_sys_tmp3809 = (w_sys_tmp3810 + r_run_k_29);
	assign w_sys_tmp3810 = 32'sh00001447;
	assign w_sys_tmp3821 = (w_sys_tmp3822 + r_run_k_29);
	assign w_sys_tmp3822 = 32'sh000014ac;
	assign w_sys_tmp3833 = (w_sys_tmp3834 + r_run_k_29);
	assign w_sys_tmp3834 = 32'sh00001511;
	assign w_sys_tmp3845 = (w_sys_tmp3846 + r_run_k_29);
	assign w_sys_tmp3846 = 32'sh00001576;
	assign w_sys_tmp3857 = (w_sys_tmp3858 + r_run_k_29);
	assign w_sys_tmp3858 = 32'sh000015db;
	assign w_sys_tmp3869 = (w_sys_tmp3870 + r_run_k_29);
	assign w_sys_tmp3870 = 32'sh00001640;
	assign w_sys_tmp3881 = (w_sys_tmp3882 + r_run_k_29);
	assign w_sys_tmp3882 = 32'sh000016a5;
	assign w_sys_tmp3893 = (w_sys_tmp3894 + r_run_k_29);
	assign w_sys_tmp3894 = 32'sh0000170a;
	assign w_sys_tmp3905 = (w_sys_tmp3906 + r_run_k_29);
	assign w_sys_tmp3906 = 32'sh0000176f;
	assign w_sys_tmp3917 = (w_sys_tmp3918 + r_run_k_29);
	assign w_sys_tmp3918 = 32'sh000017d4;
	assign w_sys_tmp3929 = (w_sys_tmp3930 + r_run_k_29);
	assign w_sys_tmp3930 = 32'sh00001839;
	assign w_sys_tmp3941 = (w_sys_tmp3942 + r_run_k_29);
	assign w_sys_tmp3942 = 32'sh0000189e;
	assign w_sys_tmp3965 = (w_sys_tmp3966 + r_run_k_29);
	assign w_sys_tmp3966 = 32'sh00001903;
	assign w_sys_tmp3977 = (w_sys_tmp3978 + r_run_k_29);
	assign w_sys_tmp3978 = 32'sh00001968;
	assign w_sys_tmp3989 = (w_sys_tmp3990 + r_run_k_29);
	assign w_sys_tmp3990 = 32'sh000019cd;
	assign w_sys_tmp4001 = (w_sys_tmp4002 + r_run_k_29);
	assign w_sys_tmp4002 = 32'sh00001a32;
	assign w_sys_tmp4013 = (w_sys_tmp4014 + r_run_k_29);
	assign w_sys_tmp4014 = 32'sh00001a97;
	assign w_sys_tmp4025 = (w_sys_tmp4026 + r_run_k_29);
	assign w_sys_tmp4026 = 32'sh00001afc;
	assign w_sys_tmp4037 = (w_sys_tmp4038 + r_run_k_29);
	assign w_sys_tmp4038 = 32'sh00001b61;
	assign w_sys_tmp4049 = (w_sys_tmp4050 + r_run_k_29);
	assign w_sys_tmp4050 = 32'sh00001bc6;
	assign w_sys_tmp4061 = (w_sys_tmp4062 + r_run_k_29);
	assign w_sys_tmp4062 = 32'sh00001c2b;
	assign w_sys_tmp4073 = (w_sys_tmp4074 + r_run_k_29);
	assign w_sys_tmp4074 = 32'sh00001c90;
	assign w_sys_tmp4085 = (w_sys_tmp4086 + r_run_k_29);
	assign w_sys_tmp4086 = 32'sh00001cf5;
	assign w_sys_tmp4097 = (w_sys_tmp4098 + r_run_k_29);
	assign w_sys_tmp4098 = 32'sh00001d5a;
	assign w_sys_tmp4109 = (w_sys_tmp4110 + r_run_k_29);
	assign w_sys_tmp4110 = 32'sh00001dbf;
	assign w_sys_tmp4121 = (w_sys_tmp4122 + r_run_k_29);
	assign w_sys_tmp4122 = 32'sh00001e24;
	assign w_sys_tmp4133 = (w_sys_tmp4134 + r_run_k_29);
	assign w_sys_tmp4134 = 32'sh00001e89;
	assign w_sys_tmp4145 = (w_sys_tmp4146 + r_run_k_29);
	assign w_sys_tmp4146 = 32'sh00001eee;
	assign w_sys_tmp4157 = (w_sys_tmp4158 + r_run_k_29);
	assign w_sys_tmp4158 = 32'sh00001f53;
	assign w_sys_tmp4169 = (w_sys_tmp4170 + r_run_k_29);
	assign w_sys_tmp4170 = 32'sh00001fb8;
	assign w_sys_tmp4181 = (w_sys_tmp4182 + r_run_k_29);
	assign w_sys_tmp4182 = 32'sh0000201d;
	assign w_sys_tmp4193 = (w_sys_tmp4194 + r_run_k_29);
	assign w_sys_tmp4194 = 32'sh00002082;
	assign w_sys_tmp4229 = (w_sys_tmp4230 + r_run_k_29);
	assign w_sys_tmp4230 = 32'sh000020e7;
	assign w_sys_tmp4241 = (w_sys_tmp4242 + r_run_k_29);
	assign w_sys_tmp4242 = 32'sh000c5dcc;
	assign w_sys_tmp4253 = (w_sys_tmp4254 + r_run_k_29);
	assign w_sys_tmp4254 = 32'sh000021b1;
	assign w_sys_tmp4265 = (w_sys_tmp4266 + r_run_k_29);
	assign w_sys_tmp4266 = 32'sh00002216;
	assign w_sys_tmp4277 = (w_sys_tmp4278 + r_run_k_29);
	assign w_sys_tmp4278 = 32'sh0000227b;
	assign w_sys_tmp4289 = (w_sys_tmp4290 + r_run_k_29);
	assign w_sys_tmp4290 = 32'sh000022e0;
	assign w_sys_tmp4301 = (w_sys_tmp4302 + r_run_k_29);
	assign w_sys_tmp4302 = 32'sh00002345;
	assign w_sys_tmp4313 = (w_sys_tmp4314 + r_run_k_29);
	assign w_sys_tmp4314 = 32'sh000023aa;
	assign w_sys_tmp4325 = (w_sys_tmp4326 + r_run_k_29);
	assign w_sys_tmp4326 = 32'sh0000240f;
	assign w_sys_tmp4337 = (w_sys_tmp4338 + r_run_k_29);
	assign w_sys_tmp4338 = 32'sh00002474;
	assign w_sys_tmp4349 = (w_sys_tmp4350 + r_run_k_29);
	assign w_sys_tmp4350 = 32'sh000024d9;
	assign w_sys_tmp4361 = (w_sys_tmp4362 + r_run_k_29);
	assign w_sys_tmp4362 = 32'sh0000253e;
	assign w_sys_tmp4373 = (w_sys_tmp4374 + r_run_k_29);
	assign w_sys_tmp4374 = 32'sh000025a3;
	assign w_sys_tmp4385 = (w_sys_tmp4386 + r_run_k_29);
	assign w_sys_tmp4386 = 32'sh00002608;
	assign w_sys_tmp4397 = (w_sys_tmp4398 + r_run_k_29);
	assign w_sys_tmp4398 = 32'sh0000266d;
	assign w_sys_tmp4409 = (w_sys_tmp4410 + r_run_k_29);
	assign w_sys_tmp4410 = 32'sh000026d2;
	assign w_sys_tmp4421 = (w_sys_tmp4422 + r_run_k_29);
	assign w_sys_tmp4422 = 32'sh00002737;
	assign w_sys_tmp4433 = (w_sys_tmp4434 + r_run_k_29);
	assign w_sys_tmp4434 = 32'sh0000279c;
	assign w_sys_tmp4445 = (w_sys_tmp4446 + r_run_k_29);
	assign w_sys_tmp4446 = 32'sh00002801;
	assign w_sys_tmp4457 = (w_sys_tmp4458 + r_run_k_29);
	assign w_sys_tmp4458 = 32'sh000000a1;
	assign w_sys_tmp4469 = (w_sys_tmp4470 + r_run_k_29);
	assign w_sys_tmp4470 = 32'sh00000106;
	assign w_sys_tmp4481 = (w_sys_tmp4482 + r_run_k_29);
	assign w_sys_tmp4482 = 32'sh0000016b;
	assign w_sys_tmp4493 = (w_sys_tmp4494 + r_run_k_29);
	assign w_sys_tmp4494 = 32'sh000001d0;
	assign w_sys_tmp4505 = (w_sys_tmp4506 + r_run_k_29);
	assign w_sys_tmp4506 = 32'sh00000235;
	assign w_sys_tmp4517 = (w_sys_tmp4518 + r_run_k_29);
	assign w_sys_tmp4518 = 32'sh0000029a;
	assign w_sys_tmp4529 = (w_sys_tmp4530 + r_run_k_29);
	assign w_sys_tmp4530 = 32'sh000002ff;
	assign w_sys_tmp4541 = (w_sys_tmp4542 + r_run_k_29);
	assign w_sys_tmp4542 = 32'sh00000364;
	assign w_sys_tmp4553 = (w_sys_tmp4554 + r_run_k_29);
	assign w_sys_tmp4554 = 32'sh000003c9;
	assign w_sys_tmp4565 = (w_sys_tmp4566 + r_run_k_29);
	assign w_sys_tmp4566 = 32'sh0000042e;
	assign w_sys_tmp4577 = (w_sys_tmp4578 + r_run_k_29);
	assign w_sys_tmp4578 = 32'sh00000493;
	assign w_sys_tmp4589 = (w_sys_tmp4590 + r_run_k_29);
	assign w_sys_tmp4590 = 32'sh000004f8;
	assign w_sys_tmp4601 = (w_sys_tmp4602 + r_run_k_29);
	assign w_sys_tmp4602 = 32'sh0000055d;
	assign w_sys_tmp4613 = (w_sys_tmp4614 + r_run_k_29);
	assign w_sys_tmp4614 = 32'sh000005c2;
	assign w_sys_tmp4625 = (w_sys_tmp4626 + r_run_k_29);
	assign w_sys_tmp4626 = 32'sh00000627;
	assign w_sys_tmp4637 = (w_sys_tmp4638 + r_run_k_29);
	assign w_sys_tmp4638 = 32'sh0000068c;
	assign w_sys_tmp4649 = (w_sys_tmp4650 + r_run_k_29);
	assign w_sys_tmp4650 = 32'sh000006f1;
	assign w_sys_tmp4661 = (w_sys_tmp4662 + r_run_k_29);
	assign w_sys_tmp4662 = 32'sh00000756;
	assign w_sys_tmp4673 = (w_sys_tmp4674 + r_run_k_29);
	assign w_sys_tmp4674 = 32'sh000007bb;
	assign w_sys_tmp4685 = (w_sys_tmp4686 + r_run_k_29);
	assign w_sys_tmp4686 = 32'sh00000820;
	assign w_sys_tmp4697 = (w_sys_tmp4698 + r_run_k_29);
	assign w_sys_tmp4698 = 32'sh00000885;
	assign w_sys_tmp4721 = (w_sys_tmp4722 + r_run_k_29);
	assign w_sys_tmp4722 = 32'sh000008ea;
	assign w_sys_tmp4733 = (w_sys_tmp4734 + r_run_k_29);
	assign w_sys_tmp4734 = 32'sh0000094f;
	assign w_sys_tmp4745 = (w_sys_tmp4746 + r_run_k_29);
	assign w_sys_tmp4746 = 32'sh000009b4;
	assign w_sys_tmp4757 = (w_sys_tmp4758 + r_run_k_29);
	assign w_sys_tmp4758 = 32'sh00000a19;
	assign w_sys_tmp4769 = (w_sys_tmp4770 + r_run_k_29);
	assign w_sys_tmp4770 = 32'sh00000a7e;
	assign w_sys_tmp4781 = (w_sys_tmp4782 + r_run_k_29);
	assign w_sys_tmp4782 = 32'sh00000ae3;
	assign w_sys_tmp4793 = (w_sys_tmp4794 + r_run_k_29);
	assign w_sys_tmp4794 = 32'sh00000b48;
	assign w_sys_tmp4805 = (w_sys_tmp4806 + r_run_k_29);
	assign w_sys_tmp4806 = 32'sh00000bad;
	assign w_sys_tmp4817 = (w_sys_tmp4818 + r_run_k_29);
	assign w_sys_tmp4818 = 32'sh00000c12;
	assign w_sys_tmp4829 = (w_sys_tmp4830 + r_run_k_29);
	assign w_sys_tmp4830 = 32'sh00000c77;
	assign w_sys_tmp4841 = (w_sys_tmp4842 + r_run_k_29);
	assign w_sys_tmp4842 = 32'sh00000cdc;
	assign w_sys_tmp4853 = (w_sys_tmp4854 + r_run_k_29);
	assign w_sys_tmp4854 = 32'sh00000d41;
	assign w_sys_tmp4865 = (w_sys_tmp4866 + r_run_k_29);
	assign w_sys_tmp4866 = 32'sh00000da6;
	assign w_sys_tmp4877 = (w_sys_tmp4878 + r_run_k_29);
	assign w_sys_tmp4878 = 32'sh00000e0b;
	assign w_sys_tmp4889 = (w_sys_tmp4890 + r_run_k_29);
	assign w_sys_tmp4890 = 32'sh00000e70;
	assign w_sys_tmp4901 = (w_sys_tmp4902 + r_run_k_29);
	assign w_sys_tmp4902 = 32'sh00000ed5;
	assign w_sys_tmp4913 = (w_sys_tmp4914 + r_run_k_29);
	assign w_sys_tmp4914 = 32'sh00000f3a;
	assign w_sys_tmp4925 = (w_sys_tmp4926 + r_run_k_29);
	assign w_sys_tmp4926 = 32'sh00000f9f;
	assign w_sys_tmp4937 = (w_sys_tmp4938 + r_run_k_29);
	assign w_sys_tmp4938 = 32'sh00001004;
	assign w_sys_tmp4949 = (w_sys_tmp4950 + r_run_k_29);
	assign w_sys_tmp4950 = 32'sh00001069;
	assign w_sys_tmp4961 = (w_sys_tmp4962 + r_run_k_29);
	assign w_sys_tmp4962 = 32'sh000010ce;
	assign w_sys_tmp4997 = (w_sys_tmp4998 + r_run_k_29);
	assign w_sys_tmp4998 = 32'sh00001133;
	assign w_sys_tmp5009 = (w_sys_tmp5010 + r_run_k_29);
	assign w_sys_tmp5010 = 32'sh00001198;
	assign w_sys_tmp5021 = (w_sys_tmp5022 + r_run_k_29);
	assign w_sys_tmp5022 = 32'sh000011fd;
	assign w_sys_tmp5033 = (w_sys_tmp5034 + r_run_k_29);
	assign w_sys_tmp5034 = 32'sh00001262;
	assign w_sys_tmp5045 = (w_sys_tmp5046 + r_run_k_29);
	assign w_sys_tmp5046 = 32'sh000012c7;
	assign w_sys_tmp5057 = (w_sys_tmp5058 + r_run_k_29);
	assign w_sys_tmp5058 = 32'sh000196ac;
	assign w_sys_tmp5069 = (w_sys_tmp5070 + r_run_k_29);
	assign w_sys_tmp5070 = 32'sh00001391;
	assign w_sys_tmp5081 = (w_sys_tmp5082 + r_run_k_29);
	assign w_sys_tmp5082 = 32'sh000013f6;
	assign w_sys_tmp5093 = (w_sys_tmp5094 + r_run_k_29);
	assign w_sys_tmp5094 = 32'sh0000145b;
	assign w_sys_tmp5105 = (w_sys_tmp5106 + r_run_k_29);
	assign w_sys_tmp5106 = 32'sh000014c0;
	assign w_sys_tmp5117 = (w_sys_tmp5118 + r_run_k_29);
	assign w_sys_tmp5118 = 32'sh00001525;
	assign w_sys_tmp5129 = (w_sys_tmp5130 + r_run_k_29);
	assign w_sys_tmp5130 = 32'sh0000158a;
	assign w_sys_tmp5141 = (w_sys_tmp5142 + r_run_k_29);
	assign w_sys_tmp5142 = 32'sh000015ef;
	assign w_sys_tmp5153 = (w_sys_tmp5154 + r_run_k_29);
	assign w_sys_tmp5154 = 32'sh00001654;
	assign w_sys_tmp5165 = (w_sys_tmp5166 + r_run_k_29);
	assign w_sys_tmp5166 = 32'sh000016b9;
	assign w_sys_tmp5177 = (w_sys_tmp5178 + r_run_k_29);
	assign w_sys_tmp5178 = 32'sh0000171e;
	assign w_sys_tmp5189 = (w_sys_tmp5190 + r_run_k_29);
	assign w_sys_tmp5190 = 32'sh00001783;
	assign w_sys_tmp5201 = (w_sys_tmp5202 + r_run_k_29);
	assign w_sys_tmp5202 = 32'sh000017e8;
	assign w_sys_tmp5213 = (w_sys_tmp5214 + r_run_k_29);
	assign w_sys_tmp5214 = 32'sh0000184d;
	assign w_sys_tmp5225 = (w_sys_tmp5226 + r_run_k_29);
	assign w_sys_tmp5226 = 32'sh000018b2;
	assign w_sys_tmp5261 = (w_sys_tmp5262 + r_run_k_29);
	assign w_sys_tmp5262 = 32'sh00001917;
	assign w_sys_tmp5273 = (w_sys_tmp5274 + r_run_k_29);
	assign w_sys_tmp5274 = 32'sh0000197c;
	assign w_sys_tmp5285 = (w_sys_tmp5286 + r_run_k_29);
	assign w_sys_tmp5286 = 32'sh000019e1;
	assign w_sys_tmp5297 = (w_sys_tmp5298 + r_run_k_29);
	assign w_sys_tmp5298 = 32'sh00001a46;
	assign w_sys_tmp5309 = (w_sys_tmp5310 + r_run_k_29);
	assign w_sys_tmp5310 = 32'sh00001aab;
	assign w_sys_tmp5321 = (w_sys_tmp5322 + r_run_k_29);
	assign w_sys_tmp5322 = 32'sh00001b10;
	assign w_sys_tmp5333 = (w_sys_tmp5334 + r_run_k_29);
	assign w_sys_tmp5334 = 32'sh00001b75;
	assign w_sys_tmp5345 = (w_sys_tmp5346 + r_run_k_29);
	assign w_sys_tmp5346 = 32'sh00001bda;
	assign w_sys_tmp5357 = (w_sys_tmp5358 + r_run_k_29);
	assign w_sys_tmp5358 = 32'sh00001c3f;
	assign w_sys_tmp5369 = (w_sys_tmp5370 + r_run_k_29);
	assign w_sys_tmp5370 = 32'sh00001ca4;
	assign w_sys_tmp5381 = (w_sys_tmp5382 + r_run_k_29);
	assign w_sys_tmp5382 = 32'sh00001d09;
	assign w_sys_tmp5393 = (w_sys_tmp5394 + r_run_k_29);
	assign w_sys_tmp5394 = 32'sh00001d6e;
	assign w_sys_tmp5405 = (w_sys_tmp5406 + r_run_k_29);
	assign w_sys_tmp5406 = 32'sh00001dd3;
	assign w_sys_tmp5417 = (w_sys_tmp5418 + r_run_k_29);
	assign w_sys_tmp5418 = 32'sh00001e38;
	assign w_sys_tmp5429 = (w_sys_tmp5430 + r_run_k_29);
	assign w_sys_tmp5430 = 32'sh00001e9d;
	assign w_sys_tmp5441 = (w_sys_tmp5442 + r_run_k_29);
	assign w_sys_tmp5442 = 32'sh00001f02;
	assign w_sys_tmp5453 = (w_sys_tmp5454 + r_run_k_29);
	assign w_sys_tmp5454 = 32'sh00001f67;
	assign w_sys_tmp5465 = (w_sys_tmp5466 + r_run_k_29);
	assign w_sys_tmp5466 = 32'sh00001fcc;
	assign w_sys_tmp5477 = (w_sys_tmp5478 + r_run_k_29);
	assign w_sys_tmp5478 = 32'sh00002031;
	assign w_sys_tmp5489 = (w_sys_tmp5490 + r_run_k_29);
	assign w_sys_tmp5490 = 32'sh00002096;
	assign w_sys_tmp5525 = (w_sys_tmp5526 + r_run_k_29);
	assign w_sys_tmp5526 = 32'sh000020fb;
	assign w_sys_tmp5537 = (w_sys_tmp5538 + r_run_k_29);
	assign w_sys_tmp5538 = 32'sh000c5de0;
	assign w_sys_tmp5549 = (w_sys_tmp5550 + r_run_k_29);
	assign w_sys_tmp5550 = 32'sh000021c5;
	assign w_sys_tmp5561 = (w_sys_tmp5562 + r_run_k_29);
	assign w_sys_tmp5562 = 32'sh0000222a;
	assign w_sys_tmp5573 = (w_sys_tmp5574 + r_run_k_29);
	assign w_sys_tmp5574 = 32'sh0000228f;
	assign w_sys_tmp5585 = (w_sys_tmp5586 + r_run_k_29);
	assign w_sys_tmp5586 = 32'sh000022f4;
	assign w_sys_tmp5597 = (w_sys_tmp5598 + r_run_k_29);
	assign w_sys_tmp5598 = 32'sh00002359;
	assign w_sys_tmp5609 = (w_sys_tmp5610 + r_run_k_29);
	assign w_sys_tmp5610 = 32'sh000023be;
	assign w_sys_tmp5621 = (w_sys_tmp5622 + r_run_k_29);
	assign w_sys_tmp5622 = 32'sh00002423;
	assign w_sys_tmp5633 = (w_sys_tmp5634 + r_run_k_29);
	assign w_sys_tmp5634 = 32'sh00002488;
	assign w_sys_tmp5645 = (w_sys_tmp5646 + r_run_k_29);
	assign w_sys_tmp5646 = 32'sh000024ed;
	assign w_sys_tmp5657 = (w_sys_tmp5658 + r_run_k_29);
	assign w_sys_tmp5658 = 32'sh00002552;
	assign w_sys_tmp5669 = (w_sys_tmp5670 + r_run_k_29);
	assign w_sys_tmp5670 = 32'sh000025b7;
	assign w_sys_tmp5681 = (w_sys_tmp5682 + r_run_k_29);
	assign w_sys_tmp5682 = 32'sh0000261c;
	assign w_sys_tmp5693 = (w_sys_tmp5694 + r_run_k_29);
	assign w_sys_tmp5694 = 32'sh00002681;
	assign w_sys_tmp5705 = (w_sys_tmp5706 + r_run_k_29);
	assign w_sys_tmp5706 = 32'sh000026e6;
	assign w_sys_tmp5717 = (w_sys_tmp5718 + r_run_k_29);
	assign w_sys_tmp5718 = 32'sh0000274b;
	assign w_sys_tmp5729 = (w_sys_tmp5730 + r_run_k_29);
	assign w_sys_tmp5730 = 32'sh000027b0;
	assign w_sys_tmp5741 = (w_sys_tmp5742 + r_run_k_29);
	assign w_sys_tmp5742 = 32'sh00002815;
	assign w_sys_tmp5752 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp5753 = 32'sh00000051;
	assign w_sys_tmp5754 = ( !w_sys_tmp5755 );
	assign w_sys_tmp5755 = (w_sys_tmp5756 < r_run_k_29);
	assign w_sys_tmp5756 = 32'sh00000065;
	assign w_sys_tmp5759 = (w_sys_tmp5760 + r_run_k_29);
	assign w_sys_tmp5760 = 32'sh00000065;
	assign w_sys_tmp5761 = w_fld_U_2_dataout_1;
	assign w_sys_tmp5767 = w_fld_V_3_dataout_1;
	assign w_sys_tmp5771 = (w_sys_tmp5772 + r_run_k_29);
	assign w_sys_tmp5772 = 32'sh000000ca;
	assign w_sys_tmp5783 = (w_sys_tmp5784 + r_run_k_29);
	assign w_sys_tmp5784 = 32'sh0000012f;
	assign w_sys_tmp5795 = (w_sys_tmp5796 + r_run_k_29);
	assign w_sys_tmp5796 = 32'sh00000194;
	assign w_sys_tmp5807 = (w_sys_tmp5808 + r_run_k_29);
	assign w_sys_tmp5808 = 32'sh000001f9;
	assign w_sys_tmp5819 = (w_sys_tmp5820 + r_run_k_29);
	assign w_sys_tmp5820 = 32'sh0000025e;
	assign w_sys_tmp5831 = (w_sys_tmp5832 + r_run_k_29);
	assign w_sys_tmp5832 = 32'sh000002c3;
	assign w_sys_tmp5843 = (w_sys_tmp5844 + r_run_k_29);
	assign w_sys_tmp5844 = 32'sh00000328;
	assign w_sys_tmp5855 = (w_sys_tmp5856 + r_run_k_29);
	assign w_sys_tmp5856 = 32'sh0000038d;
	assign w_sys_tmp5867 = (w_sys_tmp5868 + r_run_k_29);
	assign w_sys_tmp5868 = 32'sh000003f2;
	assign w_sys_tmp5879 = (w_sys_tmp5880 + r_run_k_29);
	assign w_sys_tmp5880 = 32'sh00000457;
	assign w_sys_tmp5891 = (w_sys_tmp5892 + r_run_k_29);
	assign w_sys_tmp5892 = 32'sh000004bc;
	assign w_sys_tmp5903 = (w_sys_tmp5904 + r_run_k_29);
	assign w_sys_tmp5904 = 32'sh00000521;
	assign w_sys_tmp5915 = (w_sys_tmp5916 + r_run_k_29);
	assign w_sys_tmp5916 = 32'sh00000586;
	assign w_sys_tmp5927 = (w_sys_tmp5928 + r_run_k_29);
	assign w_sys_tmp5928 = 32'sh000005eb;
	assign w_sys_tmp5939 = (w_sys_tmp5940 + r_run_k_29);
	assign w_sys_tmp5940 = 32'sh00000650;
	assign w_sys_tmp5951 = (w_sys_tmp5952 + r_run_k_29);
	assign w_sys_tmp5952 = 32'sh000006b5;
	assign w_sys_tmp5963 = (w_sys_tmp5964 + r_run_k_29);
	assign w_sys_tmp5964 = 32'sh0000071a;
	assign w_sys_tmp5975 = (w_sys_tmp5976 + r_run_k_29);
	assign w_sys_tmp5976 = 32'sh0000077f;
	assign w_sys_tmp5987 = (w_sys_tmp5988 + r_run_k_29);
	assign w_sys_tmp5988 = 32'sh000007e4;
	assign w_sys_tmp5999 = (w_sys_tmp6000 + r_run_k_29);
	assign w_sys_tmp6000 = 32'sh00000849;
	assign w_sys_tmp6023 = (w_sys_tmp6024 + r_run_k_29);
	assign w_sys_tmp6024 = 32'sh000008ae;
	assign w_sys_tmp6035 = (w_sys_tmp6036 + r_run_k_29);
	assign w_sys_tmp6036 = 32'sh00000913;
	assign w_sys_tmp6047 = (w_sys_tmp6048 + r_run_k_29);
	assign w_sys_tmp6048 = 32'sh00000978;
	assign w_sys_tmp6059 = (w_sys_tmp6060 + r_run_k_29);
	assign w_sys_tmp6060 = 32'sh000009dd;
	assign w_sys_tmp6071 = (w_sys_tmp6072 + r_run_k_29);
	assign w_sys_tmp6072 = 32'sh00000a42;
	assign w_sys_tmp6083 = (w_sys_tmp6084 + r_run_k_29);
	assign w_sys_tmp6084 = 32'sh00000aa7;
	assign w_sys_tmp6095 = (w_sys_tmp6096 + r_run_k_29);
	assign w_sys_tmp6096 = 32'sh00000b0c;
	assign w_sys_tmp6107 = (w_sys_tmp6108 + r_run_k_29);
	assign w_sys_tmp6108 = 32'sh00000b71;
	assign w_sys_tmp6119 = (w_sys_tmp6120 + r_run_k_29);
	assign w_sys_tmp6120 = 32'sh00000bd6;
	assign w_sys_tmp6131 = (w_sys_tmp6132 + r_run_k_29);
	assign w_sys_tmp6132 = 32'sh00000c3b;
	assign w_sys_tmp6143 = (w_sys_tmp6144 + r_run_k_29);
	assign w_sys_tmp6144 = 32'sh00000ca0;
	assign w_sys_tmp6155 = (w_sys_tmp6156 + r_run_k_29);
	assign w_sys_tmp6156 = 32'sh00000d05;
	assign w_sys_tmp6167 = (w_sys_tmp6168 + r_run_k_29);
	assign w_sys_tmp6168 = 32'sh00000d6a;
	assign w_sys_tmp6179 = (w_sys_tmp6180 + r_run_k_29);
	assign w_sys_tmp6180 = 32'sh00000dcf;
	assign w_sys_tmp6191 = (w_sys_tmp6192 + r_run_k_29);
	assign w_sys_tmp6192 = 32'sh00000e34;
	assign w_sys_tmp6203 = (w_sys_tmp6204 + r_run_k_29);
	assign w_sys_tmp6204 = 32'sh00000e99;
	assign w_sys_tmp6215 = (w_sys_tmp6216 + r_run_k_29);
	assign w_sys_tmp6216 = 32'sh00000efe;
	assign w_sys_tmp6227 = (w_sys_tmp6228 + r_run_k_29);
	assign w_sys_tmp6228 = 32'sh00000f63;
	assign w_sys_tmp6239 = (w_sys_tmp6240 + r_run_k_29);
	assign w_sys_tmp6240 = 32'sh00000fc8;
	assign w_sys_tmp6251 = (w_sys_tmp6252 + r_run_k_29);
	assign w_sys_tmp6252 = 32'sh0000102d;
	assign w_sys_tmp6263 = (w_sys_tmp6264 + r_run_k_29);
	assign w_sys_tmp6264 = 32'sh00001092;
	assign w_sys_tmp6299 = (w_sys_tmp6300 + r_run_k_29);
	assign w_sys_tmp6300 = 32'sh000010f7;
	assign w_sys_tmp6311 = (w_sys_tmp6312 + r_run_k_29);
	assign w_sys_tmp6312 = 32'sh0000115c;
	assign w_sys_tmp6323 = (w_sys_tmp6324 + r_run_k_29);
	assign w_sys_tmp6324 = 32'sh000011c1;
	assign w_sys_tmp6335 = (w_sys_tmp6336 + r_run_k_29);
	assign w_sys_tmp6336 = 32'sh00001226;
	assign w_sys_tmp6347 = (w_sys_tmp6348 + r_run_k_29);
	assign w_sys_tmp6348 = 32'sh0000128b;
	assign w_sys_tmp6359 = (w_sys_tmp6360 + r_run_k_29);
	assign w_sys_tmp6360 = 32'sh00019670;
	assign w_sys_tmp6371 = (w_sys_tmp6372 + r_run_k_29);
	assign w_sys_tmp6372 = 32'sh00001355;
	assign w_sys_tmp6383 = (w_sys_tmp6384 + r_run_k_29);
	assign w_sys_tmp6384 = 32'sh000013ba;
	assign w_sys_tmp6395 = (w_sys_tmp6396 + r_run_k_29);
	assign w_sys_tmp6396 = 32'sh0000141f;
	assign w_sys_tmp6407 = (w_sys_tmp6408 + r_run_k_29);
	assign w_sys_tmp6408 = 32'sh00001484;
	assign w_sys_tmp6419 = (w_sys_tmp6420 + r_run_k_29);
	assign w_sys_tmp6420 = 32'sh000014e9;
	assign w_sys_tmp6431 = (w_sys_tmp6432 + r_run_k_29);
	assign w_sys_tmp6432 = 32'sh0000154e;
	assign w_sys_tmp6443 = (w_sys_tmp6444 + r_run_k_29);
	assign w_sys_tmp6444 = 32'sh000015b3;
	assign w_sys_tmp6455 = (w_sys_tmp6456 + r_run_k_29);
	assign w_sys_tmp6456 = 32'sh00001618;
	assign w_sys_tmp6467 = (w_sys_tmp6468 + r_run_k_29);
	assign w_sys_tmp6468 = 32'sh0000167d;
	assign w_sys_tmp6479 = (w_sys_tmp6480 + r_run_k_29);
	assign w_sys_tmp6480 = 32'sh000016e2;
	assign w_sys_tmp6491 = (w_sys_tmp6492 + r_run_k_29);
	assign w_sys_tmp6492 = 32'sh00001747;
	assign w_sys_tmp6503 = (w_sys_tmp6504 + r_run_k_29);
	assign w_sys_tmp6504 = 32'sh000017ac;
	assign w_sys_tmp6515 = (w_sys_tmp6516 + r_run_k_29);
	assign w_sys_tmp6516 = 32'sh00001811;
	assign w_sys_tmp6527 = (w_sys_tmp6528 + r_run_k_29);
	assign w_sys_tmp6528 = 32'sh00001876;
	assign w_sys_tmp6563 = (w_sys_tmp6564 + r_run_k_29);
	assign w_sys_tmp6564 = 32'sh000018db;
	assign w_sys_tmp6575 = (w_sys_tmp6576 + r_run_k_29);
	assign w_sys_tmp6576 = 32'sh00001940;
	assign w_sys_tmp6587 = (w_sys_tmp6588 + r_run_k_29);
	assign w_sys_tmp6588 = 32'sh000019a5;
	assign w_sys_tmp6599 = (w_sys_tmp6600 + r_run_k_29);
	assign w_sys_tmp6600 = 32'sh00001a0a;
	assign w_sys_tmp6611 = (w_sys_tmp6612 + r_run_k_29);
	assign w_sys_tmp6612 = 32'sh00001a6f;
	assign w_sys_tmp6623 = (w_sys_tmp6624 + r_run_k_29);
	assign w_sys_tmp6624 = 32'sh00001ad4;
	assign w_sys_tmp6635 = (w_sys_tmp6636 + r_run_k_29);
	assign w_sys_tmp6636 = 32'sh00001b39;
	assign w_sys_tmp6647 = (w_sys_tmp6648 + r_run_k_29);
	assign w_sys_tmp6648 = 32'sh00001b9e;
	assign w_sys_tmp6659 = (w_sys_tmp6660 + r_run_k_29);
	assign w_sys_tmp6660 = 32'sh00001c03;
	assign w_sys_tmp6671 = (w_sys_tmp6672 + r_run_k_29);
	assign w_sys_tmp6672 = 32'sh00001c68;
	assign w_sys_tmp6683 = (w_sys_tmp6684 + r_run_k_29);
	assign w_sys_tmp6684 = 32'sh00001ccd;
	assign w_sys_tmp6695 = (w_sys_tmp6696 + r_run_k_29);
	assign w_sys_tmp6696 = 32'sh00001d32;
	assign w_sys_tmp6707 = (w_sys_tmp6708 + r_run_k_29);
	assign w_sys_tmp6708 = 32'sh00001d97;
	assign w_sys_tmp6719 = (w_sys_tmp6720 + r_run_k_29);
	assign w_sys_tmp6720 = 32'sh00001dfc;
	assign w_sys_tmp6731 = (w_sys_tmp6732 + r_run_k_29);
	assign w_sys_tmp6732 = 32'sh00001e61;
	assign w_sys_tmp6743 = (w_sys_tmp6744 + r_run_k_29);
	assign w_sys_tmp6744 = 32'sh00001ec6;
	assign w_sys_tmp6755 = (w_sys_tmp6756 + r_run_k_29);
	assign w_sys_tmp6756 = 32'sh00001f2b;
	assign w_sys_tmp6767 = (w_sys_tmp6768 + r_run_k_29);
	assign w_sys_tmp6768 = 32'sh00001f90;
	assign w_sys_tmp6779 = (w_sys_tmp6780 + r_run_k_29);
	assign w_sys_tmp6780 = 32'sh00001ff5;
	assign w_sys_tmp6791 = (w_sys_tmp6792 + r_run_k_29);
	assign w_sys_tmp6792 = 32'sh0000205a;
	assign w_sys_tmp6827 = (w_sys_tmp6828 + r_run_k_29);
	assign w_sys_tmp6828 = 32'sh000020bf;
	assign w_sys_tmp6839 = (w_sys_tmp6840 + r_run_k_29);
	assign w_sys_tmp6840 = 32'sh000c5da4;
	assign w_sys_tmp6851 = (w_sys_tmp6852 + r_run_k_29);
	assign w_sys_tmp6852 = 32'sh00002189;
	assign w_sys_tmp6863 = (w_sys_tmp6864 + r_run_k_29);
	assign w_sys_tmp6864 = 32'sh000021ee;
	assign w_sys_tmp6875 = (w_sys_tmp6876 + r_run_k_29);
	assign w_sys_tmp6876 = 32'sh00002253;
	assign w_sys_tmp6887 = (w_sys_tmp6888 + r_run_k_29);
	assign w_sys_tmp6888 = 32'sh000022b8;
	assign w_sys_tmp6899 = (w_sys_tmp6900 + r_run_k_29);
	assign w_sys_tmp6900 = 32'sh0000231d;
	assign w_sys_tmp6911 = (w_sys_tmp6912 + r_run_k_29);
	assign w_sys_tmp6912 = 32'sh00002382;
	assign w_sys_tmp6923 = (w_sys_tmp6924 + r_run_k_29);
	assign w_sys_tmp6924 = 32'sh000023e7;
	assign w_sys_tmp6935 = (w_sys_tmp6936 + r_run_k_29);
	assign w_sys_tmp6936 = 32'sh0000244c;
	assign w_sys_tmp6947 = (w_sys_tmp6948 + r_run_k_29);
	assign w_sys_tmp6948 = 32'sh000024b1;
	assign w_sys_tmp6959 = (w_sys_tmp6960 + r_run_k_29);
	assign w_sys_tmp6960 = 32'sh00002516;
	assign w_sys_tmp6971 = (w_sys_tmp6972 + r_run_k_29);
	assign w_sys_tmp6972 = 32'sh0000257b;
	assign w_sys_tmp6983 = (w_sys_tmp6984 + r_run_k_29);
	assign w_sys_tmp6984 = 32'sh000025e0;
	assign w_sys_tmp6995 = (w_sys_tmp6996 + r_run_k_29);
	assign w_sys_tmp6996 = 32'sh00002645;
	assign w_sys_tmp7007 = (w_sys_tmp7008 + r_run_k_29);
	assign w_sys_tmp7008 = 32'sh000026aa;
	assign w_sys_tmp7019 = (w_sys_tmp7020 + r_run_k_29);
	assign w_sys_tmp7020 = 32'sh0000270f;
	assign w_sys_tmp7031 = (w_sys_tmp7032 + r_run_k_29);
	assign w_sys_tmp7032 = 32'sh00002774;
	assign w_sys_tmp7043 = (w_sys_tmp7044 + r_run_k_29);
	assign w_sys_tmp7044 = 32'sh000027d9;
	assign w_sys_tmp7054 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp7055 = ( !w_sys_tmp7056 );
	assign w_sys_tmp7056 = (r_run_nlast_44 < r_run_n_31);
	assign w_sys_tmp7057 = (r_run_n_31 + w_sys_intOne);
	assign w_sys_tmp7058 = ( !w_sys_tmp7059 );
	assign w_sys_tmp7059 = (r_run_my_33 < r_run_k_29);
	assign w_sys_tmp7062 = (w_sys_tmp7063 + r_run_k_29);
	assign w_sys_tmp7063 = 32'sh00000065;
	assign w_sys_tmp7064 = 32'h0;
	assign w_sys_tmp7066 = (w_sys_tmp7067 + r_run_k_29);
	assign w_sys_tmp7067 = (r_run_mx_32 * w_sys_tmp7063);
	assign w_sys_tmp7069 = w_fld_T_0_dataout_1;
	assign w_sys_tmp7070 = (w_sys_tmp7071 + r_run_k_29);
	assign w_sys_tmp7071 = (w_sys_tmp7072 * w_sys_tmp7063);
	assign w_sys_tmp7072 = (r_run_mx_32 - w_sys_intOne);
	assign w_sys_tmp7074 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp7075 = ( !w_sys_tmp7076 );
	assign w_sys_tmp7076 = (r_run_mx_32 < r_run_j_30);
	assign w_sys_tmp7079 = (w_sys_tmp7080 + w_sys_intOne);
	assign w_sys_tmp7080 = (r_run_j_30 * w_sys_tmp7081);
	assign w_sys_tmp7081 = 32'sh00000065;
	assign w_sys_tmp7082 = 32'h0;
	assign w_sys_tmp7084 = (w_sys_tmp7085 + r_run_my_33);
	assign w_sys_tmp7085 = (r_run_copy0_j_48 * w_sys_tmp7081);
	assign w_sys_tmp7088 = (r_run_copy0_j_48 + w_sys_intOne);
	assign w_sys_tmp7089 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp7318 = w_ip_DivInt_quotient_0;
	assign w_sys_tmp7319 = 32'sh00000004;
	assign w_sys_tmp7320 = ( !w_sys_tmp7321 );
	assign w_sys_tmp7321 = (w_sys_tmp7322 < r_run_j_30);
	assign w_sys_tmp7322 = w_ip_DivInt_quotient_0;
	assign w_sys_tmp7323 = 32'sh00000002;
	assign w_sys_tmp7326 = (w_sys_tmp7327 + w_sys_intOne);
	assign w_sys_tmp7327 = (r_run_j_30 * w_sys_tmp7328);
	assign w_sys_tmp7328 = 32'sh00000065;
	assign w_sys_tmp7329 = 32'h3f800000;
	assign w_sys_tmp7330 = (r_run_j_30 + w_sys_intOne);
	assign w_sys_tmp7445 = ( !w_sys_tmp7446 );
	assign w_sys_tmp7446 = (w_sys_tmp7447 < r_run_k_29);
	assign w_sys_tmp7447 = 32'sh00000016;
	assign w_sys_tmp7450 = (w_sys_tmp7451 + r_run_k_29);
	assign w_sys_tmp7451 = 32'sh00000065;
	assign w_sys_tmp7452 = w_fld_T_0_dataout_1;
	assign w_sys_tmp7456 = (w_sys_tmp7457 + r_run_k_29);
	assign w_sys_tmp7457 = 32'sh000000ca;
	assign w_sys_tmp7462 = (w_sys_tmp7463 + r_run_k_29);
	assign w_sys_tmp7463 = 32'sh0000012f;
	assign w_sys_tmp7468 = (w_sys_tmp7469 + r_run_k_29);
	assign w_sys_tmp7469 = 32'sh00000194;
	assign w_sys_tmp7474 = (w_sys_tmp7475 + r_run_k_29);
	assign w_sys_tmp7475 = 32'sh000001f9;
	assign w_sys_tmp7480 = (w_sys_tmp7481 + r_run_k_29);
	assign w_sys_tmp7481 = 32'sh0000025e;
	assign w_sys_tmp7486 = (w_sys_tmp7487 + r_run_k_29);
	assign w_sys_tmp7487 = 32'sh000002c3;
	assign w_sys_tmp7492 = (w_sys_tmp7493 + r_run_k_29);
	assign w_sys_tmp7493 = 32'sh00000328;
	assign w_sys_tmp7498 = (w_sys_tmp7499 + r_run_k_29);
	assign w_sys_tmp7499 = 32'sh0000038d;
	assign w_sys_tmp7504 = (w_sys_tmp7505 + r_run_k_29);
	assign w_sys_tmp7505 = 32'sh000003f2;
	assign w_sys_tmp7510 = (w_sys_tmp7511 + r_run_k_29);
	assign w_sys_tmp7511 = 32'sh00000457;
	assign w_sys_tmp7516 = (w_sys_tmp7517 + r_run_k_29);
	assign w_sys_tmp7517 = 32'sh000004bc;
	assign w_sys_tmp7522 = (w_sys_tmp7523 + r_run_k_29);
	assign w_sys_tmp7523 = 32'sh00000521;
	assign w_sys_tmp7528 = (w_sys_tmp7529 + r_run_k_29);
	assign w_sys_tmp7529 = 32'sh00000586;
	assign w_sys_tmp7534 = (w_sys_tmp7535 + r_run_k_29);
	assign w_sys_tmp7535 = 32'sh000005eb;
	assign w_sys_tmp7540 = (w_sys_tmp7541 + r_run_k_29);
	assign w_sys_tmp7541 = 32'sh00000650;
	assign w_sys_tmp7546 = (w_sys_tmp7547 + r_run_k_29);
	assign w_sys_tmp7547 = 32'sh000006b5;
	assign w_sys_tmp7552 = (w_sys_tmp7553 + r_run_k_29);
	assign w_sys_tmp7553 = 32'sh0000071a;
	assign w_sys_tmp7558 = (w_sys_tmp7559 + r_run_k_29);
	assign w_sys_tmp7559 = 32'sh0000077f;
	assign w_sys_tmp7564 = (w_sys_tmp7565 + r_run_k_29);
	assign w_sys_tmp7565 = 32'sh000007e4;
	assign w_sys_tmp7570 = (w_sys_tmp7571 + r_run_k_29);
	assign w_sys_tmp7571 = 32'sh00000849;
	assign w_sys_tmp7576 = (w_sys_tmp7577 + r_run_k_29);
	assign w_sys_tmp7577 = 32'sh000008ae;
	assign w_sys_tmp7594 = (w_sys_tmp7595 + r_run_k_29);
	assign w_sys_tmp7595 = 32'sh00000913;
	assign w_sys_tmp7600 = (w_sys_tmp7601 + r_run_k_29);
	assign w_sys_tmp7601 = 32'sh00000978;
	assign w_sys_tmp7606 = (w_sys_tmp7607 + r_run_k_29);
	assign w_sys_tmp7607 = 32'sh000009dd;
	assign w_sys_tmp7612 = (w_sys_tmp7613 + r_run_k_29);
	assign w_sys_tmp7613 = 32'sh00000a42;
	assign w_sys_tmp7618 = (w_sys_tmp7619 + r_run_k_29);
	assign w_sys_tmp7619 = 32'sh00000aa7;
	assign w_sys_tmp7624 = (w_sys_tmp7625 + r_run_k_29);
	assign w_sys_tmp7625 = 32'sh00000b0c;
	assign w_sys_tmp7630 = (w_sys_tmp7631 + r_run_k_29);
	assign w_sys_tmp7631 = 32'sh00000b71;
	assign w_sys_tmp7636 = (w_sys_tmp7637 + r_run_k_29);
	assign w_sys_tmp7637 = 32'sh00000bd6;
	assign w_sys_tmp7642 = (w_sys_tmp7643 + r_run_k_29);
	assign w_sys_tmp7643 = 32'sh00000c3b;
	assign w_sys_tmp7648 = (w_sys_tmp7649 + r_run_k_29);
	assign w_sys_tmp7649 = 32'sh00000ca0;
	assign w_sys_tmp7654 = (w_sys_tmp7655 + r_run_k_29);
	assign w_sys_tmp7655 = 32'sh00000d05;
	assign w_sys_tmp7660 = (w_sys_tmp7661 + r_run_k_29);
	assign w_sys_tmp7661 = 32'sh00000d6a;
	assign w_sys_tmp7666 = (w_sys_tmp7667 + r_run_k_29);
	assign w_sys_tmp7667 = 32'sh00000dcf;
	assign w_sys_tmp7672 = (w_sys_tmp7673 + r_run_k_29);
	assign w_sys_tmp7673 = 32'sh00000e34;
	assign w_sys_tmp7678 = (w_sys_tmp7679 + r_run_k_29);
	assign w_sys_tmp7679 = 32'sh00000e99;
	assign w_sys_tmp7684 = (w_sys_tmp7685 + r_run_k_29);
	assign w_sys_tmp7685 = 32'sh00000efe;
	assign w_sys_tmp7690 = (w_sys_tmp7691 + r_run_k_29);
	assign w_sys_tmp7691 = 32'sh00000f63;
	assign w_sys_tmp7696 = (w_sys_tmp7697 + r_run_k_29);
	assign w_sys_tmp7697 = 32'sh00000fc8;
	assign w_sys_tmp7702 = (w_sys_tmp7703 + r_run_k_29);
	assign w_sys_tmp7703 = 32'sh0000102d;
	assign w_sys_tmp7708 = (w_sys_tmp7709 + r_run_k_29);
	assign w_sys_tmp7709 = 32'sh00001092;
	assign w_sys_tmp7726 = (w_sys_tmp7727 + r_run_k_29);
	assign w_sys_tmp7727 = 32'sh000010f7;
	assign w_sys_tmp7732 = (w_sys_tmp7733 + r_run_k_29);
	assign w_sys_tmp7733 = 32'sh0000115c;
	assign w_sys_tmp7738 = (w_sys_tmp7739 + r_run_k_29);
	assign w_sys_tmp7739 = 32'sh000011c1;
	assign w_sys_tmp7744 = (w_sys_tmp7745 + r_run_k_29);
	assign w_sys_tmp7745 = 32'sh00001226;
	assign w_sys_tmp7750 = (w_sys_tmp7751 + r_run_k_29);
	assign w_sys_tmp7751 = 32'sh0000128b;
	assign w_sys_tmp7756 = (w_sys_tmp7757 + r_run_k_29);
	assign w_sys_tmp7757 = 32'sh00019670;
	assign w_sys_tmp7762 = (w_sys_tmp7763 + r_run_k_29);
	assign w_sys_tmp7763 = 32'sh00001355;
	assign w_sys_tmp7768 = (w_sys_tmp7769 + r_run_k_29);
	assign w_sys_tmp7769 = 32'sh000013ba;
	assign w_sys_tmp7774 = (w_sys_tmp7775 + r_run_k_29);
	assign w_sys_tmp7775 = 32'sh0000141f;
	assign w_sys_tmp7780 = (w_sys_tmp7781 + r_run_k_29);
	assign w_sys_tmp7781 = 32'sh00001484;
	assign w_sys_tmp7786 = (w_sys_tmp7787 + r_run_k_29);
	assign w_sys_tmp7787 = 32'sh000014e9;
	assign w_sys_tmp7792 = (w_sys_tmp7793 + r_run_k_29);
	assign w_sys_tmp7793 = 32'sh0000154e;
	assign w_sys_tmp7798 = (w_sys_tmp7799 + r_run_k_29);
	assign w_sys_tmp7799 = 32'sh000015b3;
	assign w_sys_tmp7804 = (w_sys_tmp7805 + r_run_k_29);
	assign w_sys_tmp7805 = 32'sh00001618;
	assign w_sys_tmp7810 = (w_sys_tmp7811 + r_run_k_29);
	assign w_sys_tmp7811 = 32'sh0000167d;
	assign w_sys_tmp7816 = (w_sys_tmp7817 + r_run_k_29);
	assign w_sys_tmp7817 = 32'sh000016e2;
	assign w_sys_tmp7822 = (w_sys_tmp7823 + r_run_k_29);
	assign w_sys_tmp7823 = 32'sh00001747;
	assign w_sys_tmp7828 = (w_sys_tmp7829 + r_run_k_29);
	assign w_sys_tmp7829 = 32'sh000017ac;
	assign w_sys_tmp7834 = (w_sys_tmp7835 + r_run_k_29);
	assign w_sys_tmp7835 = 32'sh00001811;
	assign w_sys_tmp7840 = (w_sys_tmp7841 + r_run_k_29);
	assign w_sys_tmp7841 = 32'sh00001876;
	assign w_sys_tmp7858 = (w_sys_tmp7859 + r_run_k_29);
	assign w_sys_tmp7859 = 32'sh000018db;
	assign w_sys_tmp7864 = (w_sys_tmp7865 + r_run_k_29);
	assign w_sys_tmp7865 = 32'sh00001940;
	assign w_sys_tmp7870 = (w_sys_tmp7871 + r_run_k_29);
	assign w_sys_tmp7871 = 32'sh000019a5;
	assign w_sys_tmp7876 = (w_sys_tmp7877 + r_run_k_29);
	assign w_sys_tmp7877 = 32'sh00001a0a;
	assign w_sys_tmp7882 = (w_sys_tmp7883 + r_run_k_29);
	assign w_sys_tmp7883 = 32'sh00001a6f;
	assign w_sys_tmp7888 = (w_sys_tmp7889 + r_run_k_29);
	assign w_sys_tmp7889 = 32'sh00001ad4;
	assign w_sys_tmp7894 = (w_sys_tmp7895 + r_run_k_29);
	assign w_sys_tmp7895 = 32'sh00001b39;
	assign w_sys_tmp7900 = (w_sys_tmp7901 + r_run_k_29);
	assign w_sys_tmp7901 = 32'sh00001b9e;
	assign w_sys_tmp7906 = (w_sys_tmp7907 + r_run_k_29);
	assign w_sys_tmp7907 = 32'sh00001c03;
	assign w_sys_tmp7912 = (w_sys_tmp7913 + r_run_k_29);
	assign w_sys_tmp7913 = 32'sh00001c68;
	assign w_sys_tmp7918 = (w_sys_tmp7919 + r_run_k_29);
	assign w_sys_tmp7919 = 32'sh00001ccd;
	assign w_sys_tmp7924 = (w_sys_tmp7925 + r_run_k_29);
	assign w_sys_tmp7925 = 32'sh00001d32;
	assign w_sys_tmp7930 = (w_sys_tmp7931 + r_run_k_29);
	assign w_sys_tmp7931 = 32'sh00001d97;
	assign w_sys_tmp7936 = (w_sys_tmp7937 + r_run_k_29);
	assign w_sys_tmp7937 = 32'sh00001dfc;
	assign w_sys_tmp7942 = (w_sys_tmp7943 + r_run_k_29);
	assign w_sys_tmp7943 = 32'sh00001e61;
	assign w_sys_tmp7948 = (w_sys_tmp7949 + r_run_k_29);
	assign w_sys_tmp7949 = 32'sh00001ec6;
	assign w_sys_tmp7954 = (w_sys_tmp7955 + r_run_k_29);
	assign w_sys_tmp7955 = 32'sh00001f2b;
	assign w_sys_tmp7960 = (w_sys_tmp7961 + r_run_k_29);
	assign w_sys_tmp7961 = 32'sh00001f90;
	assign w_sys_tmp7966 = (w_sys_tmp7967 + r_run_k_29);
	assign w_sys_tmp7967 = 32'sh00001ff5;
	assign w_sys_tmp7972 = (w_sys_tmp7973 + r_run_k_29);
	assign w_sys_tmp7973 = 32'sh0000205a;
	assign w_sys_tmp7990 = (w_sys_tmp7991 + r_run_k_29);
	assign w_sys_tmp7991 = 32'sh000020bf;
	assign w_sys_tmp7996 = (w_sys_tmp7997 + r_run_k_29);
	assign w_sys_tmp7997 = 32'sh000c5da4;
	assign w_sys_tmp8002 = (w_sys_tmp8003 + r_run_k_29);
	assign w_sys_tmp8003 = 32'sh00002189;
	assign w_sys_tmp8008 = (w_sys_tmp8009 + r_run_k_29);
	assign w_sys_tmp8009 = 32'sh000021ee;
	assign w_sys_tmp8014 = (w_sys_tmp8015 + r_run_k_29);
	assign w_sys_tmp8015 = 32'sh00002253;
	assign w_sys_tmp8020 = (w_sys_tmp8021 + r_run_k_29);
	assign w_sys_tmp8021 = 32'sh000022b8;
	assign w_sys_tmp8026 = (w_sys_tmp8027 + r_run_k_29);
	assign w_sys_tmp8027 = 32'sh0000231d;
	assign w_sys_tmp8032 = (w_sys_tmp8033 + r_run_k_29);
	assign w_sys_tmp8033 = 32'sh00002382;
	assign w_sys_tmp8038 = (w_sys_tmp8039 + r_run_k_29);
	assign w_sys_tmp8039 = 32'sh000023e7;
	assign w_sys_tmp8044 = (w_sys_tmp8045 + r_run_k_29);
	assign w_sys_tmp8045 = 32'sh0000244c;
	assign w_sys_tmp8050 = (w_sys_tmp8051 + r_run_k_29);
	assign w_sys_tmp8051 = 32'sh000024b1;
	assign w_sys_tmp8056 = (w_sys_tmp8057 + r_run_k_29);
	assign w_sys_tmp8057 = 32'sh00002516;
	assign w_sys_tmp8062 = (w_sys_tmp8063 + r_run_k_29);
	assign w_sys_tmp8063 = 32'sh0000257b;
	assign w_sys_tmp8068 = (w_sys_tmp8069 + r_run_k_29);
	assign w_sys_tmp8069 = 32'sh000025e0;
	assign w_sys_tmp8074 = (w_sys_tmp8075 + r_run_k_29);
	assign w_sys_tmp8075 = 32'sh00002645;
	assign w_sys_tmp8080 = (w_sys_tmp8081 + r_run_k_29);
	assign w_sys_tmp8081 = 32'sh000026aa;
	assign w_sys_tmp8086 = (w_sys_tmp8087 + r_run_k_29);
	assign w_sys_tmp8087 = 32'sh0000270f;
	assign w_sys_tmp8092 = (w_sys_tmp8093 + r_run_k_29);
	assign w_sys_tmp8093 = 32'sh00002774;
	assign w_sys_tmp8098 = (w_sys_tmp8099 + r_run_k_29);
	assign w_sys_tmp8099 = 32'sh000027d9;
	assign w_sys_tmp8104 = (w_sys_tmp8105 + r_run_k_29);
	assign w_sys_tmp8105 = 32'sh00000079;
	assign w_sys_tmp8110 = (w_sys_tmp8111 + r_run_k_29);
	assign w_sys_tmp8111 = 32'sh000000de;
	assign w_sys_tmp8116 = (w_sys_tmp8117 + r_run_k_29);
	assign w_sys_tmp8117 = 32'sh00000143;
	assign w_sys_tmp8122 = (w_sys_tmp8123 + r_run_k_29);
	assign w_sys_tmp8123 = 32'sh000001a8;
	assign w_sys_tmp8128 = (w_sys_tmp8129 + r_run_k_29);
	assign w_sys_tmp8129 = 32'sh0000020d;
	assign w_sys_tmp8134 = (w_sys_tmp8135 + r_run_k_29);
	assign w_sys_tmp8135 = 32'sh00000272;
	assign w_sys_tmp8140 = (w_sys_tmp8141 + r_run_k_29);
	assign w_sys_tmp8141 = 32'sh000002d7;
	assign w_sys_tmp8146 = (w_sys_tmp8147 + r_run_k_29);
	assign w_sys_tmp8147 = 32'sh0000033c;
	assign w_sys_tmp8152 = (w_sys_tmp8153 + r_run_k_29);
	assign w_sys_tmp8153 = 32'sh000003a1;
	assign w_sys_tmp8158 = (w_sys_tmp8159 + r_run_k_29);
	assign w_sys_tmp8159 = 32'sh00000406;
	assign w_sys_tmp8164 = (w_sys_tmp8165 + r_run_k_29);
	assign w_sys_tmp8165 = 32'sh0000046b;
	assign w_sys_tmp8170 = (w_sys_tmp8171 + r_run_k_29);
	assign w_sys_tmp8171 = 32'sh000004d0;
	assign w_sys_tmp8176 = (w_sys_tmp8177 + r_run_k_29);
	assign w_sys_tmp8177 = 32'sh00000535;
	assign w_sys_tmp8182 = (w_sys_tmp8183 + r_run_k_29);
	assign w_sys_tmp8183 = 32'sh0000059a;
	assign w_sys_tmp8188 = (w_sys_tmp8189 + r_run_k_29);
	assign w_sys_tmp8189 = 32'sh000005ff;
	assign w_sys_tmp8194 = (w_sys_tmp8195 + r_run_k_29);
	assign w_sys_tmp8195 = 32'sh00000664;
	assign w_sys_tmp8200 = (w_sys_tmp8201 + r_run_k_29);
	assign w_sys_tmp8201 = 32'sh000006c9;
	assign w_sys_tmp8206 = (w_sys_tmp8207 + r_run_k_29);
	assign w_sys_tmp8207 = 32'sh0000072e;
	assign w_sys_tmp8212 = (w_sys_tmp8213 + r_run_k_29);
	assign w_sys_tmp8213 = 32'sh00000793;
	assign w_sys_tmp8218 = (w_sys_tmp8219 + r_run_k_29);
	assign w_sys_tmp8219 = 32'sh000007f8;
	assign w_sys_tmp8224 = (w_sys_tmp8225 + r_run_k_29);
	assign w_sys_tmp8225 = 32'sh0000085d;
	assign w_sys_tmp8230 = (w_sys_tmp8231 + r_run_k_29);
	assign w_sys_tmp8231 = 32'sh000008c2;
	assign w_sys_tmp8248 = (w_sys_tmp8249 + r_run_k_29);
	assign w_sys_tmp8249 = 32'sh00000927;
	assign w_sys_tmp8254 = (w_sys_tmp8255 + r_run_k_29);
	assign w_sys_tmp8255 = 32'sh0000098c;
	assign w_sys_tmp8260 = (w_sys_tmp8261 + r_run_k_29);
	assign w_sys_tmp8261 = 32'sh000009f1;
	assign w_sys_tmp8266 = (w_sys_tmp8267 + r_run_k_29);
	assign w_sys_tmp8267 = 32'sh00000a56;
	assign w_sys_tmp8272 = (w_sys_tmp8273 + r_run_k_29);
	assign w_sys_tmp8273 = 32'sh00000abb;
	assign w_sys_tmp8278 = (w_sys_tmp8279 + r_run_k_29);
	assign w_sys_tmp8279 = 32'sh00000b20;
	assign w_sys_tmp8284 = (w_sys_tmp8285 + r_run_k_29);
	assign w_sys_tmp8285 = 32'sh00000b85;
	assign w_sys_tmp8290 = (w_sys_tmp8291 + r_run_k_29);
	assign w_sys_tmp8291 = 32'sh00000bea;
	assign w_sys_tmp8296 = (w_sys_tmp8297 + r_run_k_29);
	assign w_sys_tmp8297 = 32'sh00000c4f;
	assign w_sys_tmp8302 = (w_sys_tmp8303 + r_run_k_29);
	assign w_sys_tmp8303 = 32'sh00000cb4;
	assign w_sys_tmp8308 = (w_sys_tmp8309 + r_run_k_29);
	assign w_sys_tmp8309 = 32'sh00000d19;
	assign w_sys_tmp8314 = (w_sys_tmp8315 + r_run_k_29);
	assign w_sys_tmp8315 = 32'sh00000d7e;
	assign w_sys_tmp8320 = (w_sys_tmp8321 + r_run_k_29);
	assign w_sys_tmp8321 = 32'sh00000de3;
	assign w_sys_tmp8326 = (w_sys_tmp8327 + r_run_k_29);
	assign w_sys_tmp8327 = 32'sh00000e48;
	assign w_sys_tmp8332 = (w_sys_tmp8333 + r_run_k_29);
	assign w_sys_tmp8333 = 32'sh00000ead;
	assign w_sys_tmp8338 = (w_sys_tmp8339 + r_run_k_29);
	assign w_sys_tmp8339 = 32'sh00000f12;
	assign w_sys_tmp8344 = (w_sys_tmp8345 + r_run_k_29);
	assign w_sys_tmp8345 = 32'sh00000f77;
	assign w_sys_tmp8350 = (w_sys_tmp8351 + r_run_k_29);
	assign w_sys_tmp8351 = 32'sh00000fdc;
	assign w_sys_tmp8356 = (w_sys_tmp8357 + r_run_k_29);
	assign w_sys_tmp8357 = 32'sh00001041;
	assign w_sys_tmp8362 = (w_sys_tmp8363 + r_run_k_29);
	assign w_sys_tmp8363 = 32'sh000010a6;
	assign w_sys_tmp8380 = (w_sys_tmp8381 + r_run_k_29);
	assign w_sys_tmp8381 = 32'sh0000110b;
	assign w_sys_tmp8386 = (w_sys_tmp8387 + r_run_k_29);
	assign w_sys_tmp8387 = 32'sh00001170;
	assign w_sys_tmp8392 = (w_sys_tmp8393 + r_run_k_29);
	assign w_sys_tmp8393 = 32'sh000011d5;
	assign w_sys_tmp8398 = (w_sys_tmp8399 + r_run_k_29);
	assign w_sys_tmp8399 = 32'sh0000123a;
	assign w_sys_tmp8404 = (w_sys_tmp8405 + r_run_k_29);
	assign w_sys_tmp8405 = 32'sh0000129f;
	assign w_sys_tmp8410 = (w_sys_tmp8411 + r_run_k_29);
	assign w_sys_tmp8411 = 32'sh00019684;
	assign w_sys_tmp8416 = (w_sys_tmp8417 + r_run_k_29);
	assign w_sys_tmp8417 = 32'sh00001369;
	assign w_sys_tmp8422 = (w_sys_tmp8423 + r_run_k_29);
	assign w_sys_tmp8423 = 32'sh000013ce;
	assign w_sys_tmp8428 = (w_sys_tmp8429 + r_run_k_29);
	assign w_sys_tmp8429 = 32'sh00001433;
	assign w_sys_tmp8434 = (w_sys_tmp8435 + r_run_k_29);
	assign w_sys_tmp8435 = 32'sh00001498;
	assign w_sys_tmp8440 = (w_sys_tmp8441 + r_run_k_29);
	assign w_sys_tmp8441 = 32'sh000014fd;
	assign w_sys_tmp8446 = (w_sys_tmp8447 + r_run_k_29);
	assign w_sys_tmp8447 = 32'sh00001562;
	assign w_sys_tmp8452 = (w_sys_tmp8453 + r_run_k_29);
	assign w_sys_tmp8453 = 32'sh000015c7;
	assign w_sys_tmp8458 = (w_sys_tmp8459 + r_run_k_29);
	assign w_sys_tmp8459 = 32'sh0000162c;
	assign w_sys_tmp8464 = (w_sys_tmp8465 + r_run_k_29);
	assign w_sys_tmp8465 = 32'sh00001691;
	assign w_sys_tmp8470 = (w_sys_tmp8471 + r_run_k_29);
	assign w_sys_tmp8471 = 32'sh000016f6;
	assign w_sys_tmp8476 = (w_sys_tmp8477 + r_run_k_29);
	assign w_sys_tmp8477 = 32'sh0000175b;
	assign w_sys_tmp8482 = (w_sys_tmp8483 + r_run_k_29);
	assign w_sys_tmp8483 = 32'sh000017c0;
	assign w_sys_tmp8488 = (w_sys_tmp8489 + r_run_k_29);
	assign w_sys_tmp8489 = 32'sh00001825;
	assign w_sys_tmp8494 = (w_sys_tmp8495 + r_run_k_29);
	assign w_sys_tmp8495 = 32'sh0000188a;
	assign w_sys_tmp8512 = (w_sys_tmp8513 + r_run_k_29);
	assign w_sys_tmp8513 = 32'sh000018ef;
	assign w_sys_tmp8518 = (w_sys_tmp8519 + r_run_k_29);
	assign w_sys_tmp8519 = 32'sh00001954;
	assign w_sys_tmp8524 = (w_sys_tmp8525 + r_run_k_29);
	assign w_sys_tmp8525 = 32'sh000019b9;
	assign w_sys_tmp8530 = (w_sys_tmp8531 + r_run_k_29);
	assign w_sys_tmp8531 = 32'sh00001a1e;
	assign w_sys_tmp8536 = (w_sys_tmp8537 + r_run_k_29);
	assign w_sys_tmp8537 = 32'sh00001a83;
	assign w_sys_tmp8542 = (w_sys_tmp8543 + r_run_k_29);
	assign w_sys_tmp8543 = 32'sh00001ae8;
	assign w_sys_tmp8548 = (w_sys_tmp8549 + r_run_k_29);
	assign w_sys_tmp8549 = 32'sh00001b4d;
	assign w_sys_tmp8554 = (w_sys_tmp8555 + r_run_k_29);
	assign w_sys_tmp8555 = 32'sh00001bb2;
	assign w_sys_tmp8560 = (w_sys_tmp8561 + r_run_k_29);
	assign w_sys_tmp8561 = 32'sh00001c17;
	assign w_sys_tmp8566 = (w_sys_tmp8567 + r_run_k_29);
	assign w_sys_tmp8567 = 32'sh00001c7c;
	assign w_sys_tmp8572 = (w_sys_tmp8573 + r_run_k_29);
	assign w_sys_tmp8573 = 32'sh00001ce1;
	assign w_sys_tmp8578 = (w_sys_tmp8579 + r_run_k_29);
	assign w_sys_tmp8579 = 32'sh00001d46;
	assign w_sys_tmp8584 = (w_sys_tmp8585 + r_run_k_29);
	assign w_sys_tmp8585 = 32'sh00001dab;
	assign w_sys_tmp8590 = (w_sys_tmp8591 + r_run_k_29);
	assign w_sys_tmp8591 = 32'sh00001e10;
	assign w_sys_tmp8596 = (w_sys_tmp8597 + r_run_k_29);
	assign w_sys_tmp8597 = 32'sh00001e75;
	assign w_sys_tmp8602 = (w_sys_tmp8603 + r_run_k_29);
	assign w_sys_tmp8603 = 32'sh00001eda;
	assign w_sys_tmp8608 = (w_sys_tmp8609 + r_run_k_29);
	assign w_sys_tmp8609 = 32'sh00001f3f;
	assign w_sys_tmp8614 = (w_sys_tmp8615 + r_run_k_29);
	assign w_sys_tmp8615 = 32'sh00001fa4;
	assign w_sys_tmp8620 = (w_sys_tmp8621 + r_run_k_29);
	assign w_sys_tmp8621 = 32'sh00002009;
	assign w_sys_tmp8626 = (w_sys_tmp8627 + r_run_k_29);
	assign w_sys_tmp8627 = 32'sh0000206e;
	assign w_sys_tmp8644 = (w_sys_tmp8645 + r_run_k_29);
	assign w_sys_tmp8645 = 32'sh000020d3;
	assign w_sys_tmp8650 = (w_sys_tmp8651 + r_run_k_29);
	assign w_sys_tmp8651 = 32'sh000c5db8;
	assign w_sys_tmp8656 = (w_sys_tmp8657 + r_run_k_29);
	assign w_sys_tmp8657 = 32'sh0000219d;
	assign w_sys_tmp8662 = (w_sys_tmp8663 + r_run_k_29);
	assign w_sys_tmp8663 = 32'sh00002202;
	assign w_sys_tmp8668 = (w_sys_tmp8669 + r_run_k_29);
	assign w_sys_tmp8669 = 32'sh00002267;
	assign w_sys_tmp8674 = (w_sys_tmp8675 + r_run_k_29);
	assign w_sys_tmp8675 = 32'sh000022cc;
	assign w_sys_tmp8680 = (w_sys_tmp8681 + r_run_k_29);
	assign w_sys_tmp8681 = 32'sh00002331;
	assign w_sys_tmp8686 = (w_sys_tmp8687 + r_run_k_29);
	assign w_sys_tmp8687 = 32'sh00002396;
	assign w_sys_tmp8692 = (w_sys_tmp8693 + r_run_k_29);
	assign w_sys_tmp8693 = 32'sh000023fb;
	assign w_sys_tmp8698 = (w_sys_tmp8699 + r_run_k_29);
	assign w_sys_tmp8699 = 32'sh00002460;
	assign w_sys_tmp8704 = (w_sys_tmp8705 + r_run_k_29);
	assign w_sys_tmp8705 = 32'sh000024c5;
	assign w_sys_tmp8710 = (w_sys_tmp8711 + r_run_k_29);
	assign w_sys_tmp8711 = 32'sh0000252a;
	assign w_sys_tmp8716 = (w_sys_tmp8717 + r_run_k_29);
	assign w_sys_tmp8717 = 32'sh0000258f;
	assign w_sys_tmp8722 = (w_sys_tmp8723 + r_run_k_29);
	assign w_sys_tmp8723 = 32'sh000025f4;
	assign w_sys_tmp8728 = (w_sys_tmp8729 + r_run_k_29);
	assign w_sys_tmp8729 = 32'sh00002659;
	assign w_sys_tmp8734 = (w_sys_tmp8735 + r_run_k_29);
	assign w_sys_tmp8735 = 32'sh000026be;
	assign w_sys_tmp8740 = (w_sys_tmp8741 + r_run_k_29);
	assign w_sys_tmp8741 = 32'sh00002723;
	assign w_sys_tmp8746 = (w_sys_tmp8747 + r_run_k_29);
	assign w_sys_tmp8747 = 32'sh00002788;
	assign w_sys_tmp8752 = (w_sys_tmp8753 + r_run_k_29);
	assign w_sys_tmp8753 = 32'sh000027ed;
	assign w_sys_tmp8758 = (w_sys_tmp8759 + r_run_k_29);
	assign w_sys_tmp8759 = 32'sh0000008d;
	assign w_sys_tmp8764 = (w_sys_tmp8765 + r_run_k_29);
	assign w_sys_tmp8765 = 32'sh000000f2;
	assign w_sys_tmp8770 = (w_sys_tmp8771 + r_run_k_29);
	assign w_sys_tmp8771 = 32'sh00000157;
	assign w_sys_tmp8776 = (w_sys_tmp8777 + r_run_k_29);
	assign w_sys_tmp8777 = 32'sh000001bc;
	assign w_sys_tmp8782 = (w_sys_tmp8783 + r_run_k_29);
	assign w_sys_tmp8783 = 32'sh00000221;
	assign w_sys_tmp8788 = (w_sys_tmp8789 + r_run_k_29);
	assign w_sys_tmp8789 = 32'sh00000286;
	assign w_sys_tmp8794 = (w_sys_tmp8795 + r_run_k_29);
	assign w_sys_tmp8795 = 32'sh000002eb;
	assign w_sys_tmp8800 = (w_sys_tmp8801 + r_run_k_29);
	assign w_sys_tmp8801 = 32'sh00000350;
	assign w_sys_tmp8806 = (w_sys_tmp8807 + r_run_k_29);
	assign w_sys_tmp8807 = 32'sh000003b5;
	assign w_sys_tmp8812 = (w_sys_tmp8813 + r_run_k_29);
	assign w_sys_tmp8813 = 32'sh0000041a;
	assign w_sys_tmp8818 = (w_sys_tmp8819 + r_run_k_29);
	assign w_sys_tmp8819 = 32'sh0000047f;
	assign w_sys_tmp8824 = (w_sys_tmp8825 + r_run_k_29);
	assign w_sys_tmp8825 = 32'sh000004e4;
	assign w_sys_tmp8830 = (w_sys_tmp8831 + r_run_k_29);
	assign w_sys_tmp8831 = 32'sh00000549;
	assign w_sys_tmp8836 = (w_sys_tmp8837 + r_run_k_29);
	assign w_sys_tmp8837 = 32'sh000005ae;
	assign w_sys_tmp8842 = (w_sys_tmp8843 + r_run_k_29);
	assign w_sys_tmp8843 = 32'sh00000613;
	assign w_sys_tmp8848 = (w_sys_tmp8849 + r_run_k_29);
	assign w_sys_tmp8849 = 32'sh00000678;
	assign w_sys_tmp8854 = (w_sys_tmp8855 + r_run_k_29);
	assign w_sys_tmp8855 = 32'sh000006dd;
	assign w_sys_tmp8860 = (w_sys_tmp8861 + r_run_k_29);
	assign w_sys_tmp8861 = 32'sh00000742;
	assign w_sys_tmp8866 = (w_sys_tmp8867 + r_run_k_29);
	assign w_sys_tmp8867 = 32'sh000007a7;
	assign w_sys_tmp8872 = (w_sys_tmp8873 + r_run_k_29);
	assign w_sys_tmp8873 = 32'sh0000080c;
	assign w_sys_tmp8878 = (w_sys_tmp8879 + r_run_k_29);
	assign w_sys_tmp8879 = 32'sh00000871;
	assign w_sys_tmp8884 = (w_sys_tmp8885 + r_run_k_29);
	assign w_sys_tmp8885 = 32'sh000008d6;
	assign w_sys_tmp8902 = (w_sys_tmp8903 + r_run_k_29);
	assign w_sys_tmp8903 = 32'sh0000093b;
	assign w_sys_tmp8908 = (w_sys_tmp8909 + r_run_k_29);
	assign w_sys_tmp8909 = 32'sh000009a0;
	assign w_sys_tmp8914 = (w_sys_tmp8915 + r_run_k_29);
	assign w_sys_tmp8915 = 32'sh00000a05;
	assign w_sys_tmp8920 = (w_sys_tmp8921 + r_run_k_29);
	assign w_sys_tmp8921 = 32'sh00000a6a;
	assign w_sys_tmp8926 = (w_sys_tmp8927 + r_run_k_29);
	assign w_sys_tmp8927 = 32'sh00000acf;
	assign w_sys_tmp8932 = (w_sys_tmp8933 + r_run_k_29);
	assign w_sys_tmp8933 = 32'sh00000b34;
	assign w_sys_tmp8938 = (w_sys_tmp8939 + r_run_k_29);
	assign w_sys_tmp8939 = 32'sh00000b99;
	assign w_sys_tmp8944 = (w_sys_tmp8945 + r_run_k_29);
	assign w_sys_tmp8945 = 32'sh00000bfe;
	assign w_sys_tmp8950 = (w_sys_tmp8951 + r_run_k_29);
	assign w_sys_tmp8951 = 32'sh00000c63;
	assign w_sys_tmp8956 = (w_sys_tmp8957 + r_run_k_29);
	assign w_sys_tmp8957 = 32'sh00000cc8;
	assign w_sys_tmp8962 = (w_sys_tmp8963 + r_run_k_29);
	assign w_sys_tmp8963 = 32'sh00000d2d;
	assign w_sys_tmp8968 = (w_sys_tmp8969 + r_run_k_29);
	assign w_sys_tmp8969 = 32'sh00000d92;
	assign w_sys_tmp8974 = (w_sys_tmp8975 + r_run_k_29);
	assign w_sys_tmp8975 = 32'sh00000df7;
	assign w_sys_tmp8980 = (w_sys_tmp8981 + r_run_k_29);
	assign w_sys_tmp8981 = 32'sh00000e5c;
	assign w_sys_tmp8986 = (w_sys_tmp8987 + r_run_k_29);
	assign w_sys_tmp8987 = 32'sh00000ec1;
	assign w_sys_tmp8992 = (w_sys_tmp8993 + r_run_k_29);
	assign w_sys_tmp8993 = 32'sh00000f26;
	assign w_sys_tmp8998 = (w_sys_tmp8999 + r_run_k_29);
	assign w_sys_tmp8999 = 32'sh00000f8b;
	assign w_sys_tmp9004 = (w_sys_tmp9005 + r_run_k_29);
	assign w_sys_tmp9005 = 32'sh00000ff0;
	assign w_sys_tmp9010 = (w_sys_tmp9011 + r_run_k_29);
	assign w_sys_tmp9011 = 32'sh00001055;
	assign w_sys_tmp9016 = (w_sys_tmp9017 + r_run_k_29);
	assign w_sys_tmp9017 = 32'sh000010ba;
	assign w_sys_tmp9034 = (w_sys_tmp9035 + r_run_k_29);
	assign w_sys_tmp9035 = 32'sh0000111f;
	assign w_sys_tmp9040 = (w_sys_tmp9041 + r_run_k_29);
	assign w_sys_tmp9041 = 32'sh00001184;
	assign w_sys_tmp9046 = (w_sys_tmp9047 + r_run_k_29);
	assign w_sys_tmp9047 = 32'sh000011e9;
	assign w_sys_tmp9052 = (w_sys_tmp9053 + r_run_k_29);
	assign w_sys_tmp9053 = 32'sh0000124e;
	assign w_sys_tmp9058 = (w_sys_tmp9059 + r_run_k_29);
	assign w_sys_tmp9059 = 32'sh000012b3;
	assign w_sys_tmp9064 = (w_sys_tmp9065 + r_run_k_29);
	assign w_sys_tmp9065 = 32'sh00019698;
	assign w_sys_tmp9070 = (w_sys_tmp9071 + r_run_k_29);
	assign w_sys_tmp9071 = 32'sh0000137d;
	assign w_sys_tmp9076 = (w_sys_tmp9077 + r_run_k_29);
	assign w_sys_tmp9077 = 32'sh000013e2;
	assign w_sys_tmp9082 = (w_sys_tmp9083 + r_run_k_29);
	assign w_sys_tmp9083 = 32'sh00001447;
	assign w_sys_tmp9088 = (w_sys_tmp9089 + r_run_k_29);
	assign w_sys_tmp9089 = 32'sh000014ac;
	assign w_sys_tmp9094 = (w_sys_tmp9095 + r_run_k_29);
	assign w_sys_tmp9095 = 32'sh00001511;
	assign w_sys_tmp9100 = (w_sys_tmp9101 + r_run_k_29);
	assign w_sys_tmp9101 = 32'sh00001576;
	assign w_sys_tmp9106 = (w_sys_tmp9107 + r_run_k_29);
	assign w_sys_tmp9107 = 32'sh000015db;
	assign w_sys_tmp9112 = (w_sys_tmp9113 + r_run_k_29);
	assign w_sys_tmp9113 = 32'sh00001640;
	assign w_sys_tmp9118 = (w_sys_tmp9119 + r_run_k_29);
	assign w_sys_tmp9119 = 32'sh000016a5;
	assign w_sys_tmp9124 = (w_sys_tmp9125 + r_run_k_29);
	assign w_sys_tmp9125 = 32'sh0000170a;
	assign w_sys_tmp9130 = (w_sys_tmp9131 + r_run_k_29);
	assign w_sys_tmp9131 = 32'sh0000176f;
	assign w_sys_tmp9136 = (w_sys_tmp9137 + r_run_k_29);
	assign w_sys_tmp9137 = 32'sh000017d4;
	assign w_sys_tmp9142 = (w_sys_tmp9143 + r_run_k_29);
	assign w_sys_tmp9143 = 32'sh00001839;
	assign w_sys_tmp9148 = (w_sys_tmp9149 + r_run_k_29);
	assign w_sys_tmp9149 = 32'sh0000189e;
	assign w_sys_tmp9166 = (w_sys_tmp9167 + r_run_k_29);
	assign w_sys_tmp9167 = 32'sh00001903;
	assign w_sys_tmp9172 = (w_sys_tmp9173 + r_run_k_29);
	assign w_sys_tmp9173 = 32'sh00001968;
	assign w_sys_tmp9178 = (w_sys_tmp9179 + r_run_k_29);
	assign w_sys_tmp9179 = 32'sh000019cd;
	assign w_sys_tmp9184 = (w_sys_tmp9185 + r_run_k_29);
	assign w_sys_tmp9185 = 32'sh00001a32;
	assign w_sys_tmp9190 = (w_sys_tmp9191 + r_run_k_29);
	assign w_sys_tmp9191 = 32'sh00001a97;
	assign w_sys_tmp9196 = (w_sys_tmp9197 + r_run_k_29);
	assign w_sys_tmp9197 = 32'sh00001afc;
	assign w_sys_tmp9202 = (w_sys_tmp9203 + r_run_k_29);
	assign w_sys_tmp9203 = 32'sh00001b61;
	assign w_sys_tmp9208 = (w_sys_tmp9209 + r_run_k_29);
	assign w_sys_tmp9209 = 32'sh00001bc6;
	assign w_sys_tmp9214 = (w_sys_tmp9215 + r_run_k_29);
	assign w_sys_tmp9215 = 32'sh00001c2b;
	assign w_sys_tmp9220 = (w_sys_tmp9221 + r_run_k_29);
	assign w_sys_tmp9221 = 32'sh00001c90;
	assign w_sys_tmp9226 = (w_sys_tmp9227 + r_run_k_29);
	assign w_sys_tmp9227 = 32'sh00001cf5;
	assign w_sys_tmp9232 = (w_sys_tmp9233 + r_run_k_29);
	assign w_sys_tmp9233 = 32'sh00001d5a;
	assign w_sys_tmp9238 = (w_sys_tmp9239 + r_run_k_29);
	assign w_sys_tmp9239 = 32'sh00001dbf;
	assign w_sys_tmp9244 = (w_sys_tmp9245 + r_run_k_29);
	assign w_sys_tmp9245 = 32'sh00001e24;
	assign w_sys_tmp9250 = (w_sys_tmp9251 + r_run_k_29);
	assign w_sys_tmp9251 = 32'sh00001e89;
	assign w_sys_tmp9256 = (w_sys_tmp9257 + r_run_k_29);
	assign w_sys_tmp9257 = 32'sh00001eee;
	assign w_sys_tmp9262 = (w_sys_tmp9263 + r_run_k_29);
	assign w_sys_tmp9263 = 32'sh00001f53;
	assign w_sys_tmp9268 = (w_sys_tmp9269 + r_run_k_29);
	assign w_sys_tmp9269 = 32'sh00001fb8;
	assign w_sys_tmp9274 = (w_sys_tmp9275 + r_run_k_29);
	assign w_sys_tmp9275 = 32'sh0000201d;
	assign w_sys_tmp9280 = (w_sys_tmp9281 + r_run_k_29);
	assign w_sys_tmp9281 = 32'sh00002082;
	assign w_sys_tmp9298 = (w_sys_tmp9299 + r_run_k_29);
	assign w_sys_tmp9299 = 32'sh000020e7;
	assign w_sys_tmp9304 = (w_sys_tmp9305 + r_run_k_29);
	assign w_sys_tmp9305 = 32'sh000c5dcc;
	assign w_sys_tmp9310 = (w_sys_tmp9311 + r_run_k_29);
	assign w_sys_tmp9311 = 32'sh000021b1;
	assign w_sys_tmp9316 = (w_sys_tmp9317 + r_run_k_29);
	assign w_sys_tmp9317 = 32'sh00002216;
	assign w_sys_tmp9322 = (w_sys_tmp9323 + r_run_k_29);
	assign w_sys_tmp9323 = 32'sh0000227b;
	assign w_sys_tmp9328 = (w_sys_tmp9329 + r_run_k_29);
	assign w_sys_tmp9329 = 32'sh000022e0;
	assign w_sys_tmp9334 = (w_sys_tmp9335 + r_run_k_29);
	assign w_sys_tmp9335 = 32'sh00002345;
	assign w_sys_tmp9340 = (w_sys_tmp9341 + r_run_k_29);
	assign w_sys_tmp9341 = 32'sh000023aa;
	assign w_sys_tmp9346 = (w_sys_tmp9347 + r_run_k_29);
	assign w_sys_tmp9347 = 32'sh0000240f;
	assign w_sys_tmp9352 = (w_sys_tmp9353 + r_run_k_29);
	assign w_sys_tmp9353 = 32'sh00002474;
	assign w_sys_tmp9358 = (w_sys_tmp9359 + r_run_k_29);
	assign w_sys_tmp9359 = 32'sh000024d9;
	assign w_sys_tmp9364 = (w_sys_tmp9365 + r_run_k_29);
	assign w_sys_tmp9365 = 32'sh0000253e;
	assign w_sys_tmp9370 = (w_sys_tmp9371 + r_run_k_29);
	assign w_sys_tmp9371 = 32'sh000025a3;
	assign w_sys_tmp9376 = (w_sys_tmp9377 + r_run_k_29);
	assign w_sys_tmp9377 = 32'sh00002608;
	assign w_sys_tmp9382 = (w_sys_tmp9383 + r_run_k_29);
	assign w_sys_tmp9383 = 32'sh0000266d;
	assign w_sys_tmp9388 = (w_sys_tmp9389 + r_run_k_29);
	assign w_sys_tmp9389 = 32'sh000026d2;
	assign w_sys_tmp9394 = (w_sys_tmp9395 + r_run_k_29);
	assign w_sys_tmp9395 = 32'sh00002737;
	assign w_sys_tmp9400 = (w_sys_tmp9401 + r_run_k_29);
	assign w_sys_tmp9401 = 32'sh0000279c;
	assign w_sys_tmp9406 = (w_sys_tmp9407 + r_run_k_29);
	assign w_sys_tmp9407 = 32'sh00002801;
	assign w_sys_tmp9412 = (w_sys_tmp9413 + r_run_k_29);
	assign w_sys_tmp9413 = 32'sh000000a1;
	assign w_sys_tmp9418 = (w_sys_tmp9419 + r_run_k_29);
	assign w_sys_tmp9419 = 32'sh00000106;
	assign w_sys_tmp9424 = (w_sys_tmp9425 + r_run_k_29);
	assign w_sys_tmp9425 = 32'sh0000016b;
	assign w_sys_tmp9430 = (w_sys_tmp9431 + r_run_k_29);
	assign w_sys_tmp9431 = 32'sh000001d0;
	assign w_sys_tmp9436 = (w_sys_tmp9437 + r_run_k_29);
	assign w_sys_tmp9437 = 32'sh00000235;
	assign w_sys_tmp9442 = (w_sys_tmp9443 + r_run_k_29);
	assign w_sys_tmp9443 = 32'sh0000029a;
	assign w_sys_tmp9448 = (w_sys_tmp9449 + r_run_k_29);
	assign w_sys_tmp9449 = 32'sh000002ff;
	assign w_sys_tmp9454 = (w_sys_tmp9455 + r_run_k_29);
	assign w_sys_tmp9455 = 32'sh00000364;
	assign w_sys_tmp9460 = (w_sys_tmp9461 + r_run_k_29);
	assign w_sys_tmp9461 = 32'sh000003c9;
	assign w_sys_tmp9466 = (w_sys_tmp9467 + r_run_k_29);
	assign w_sys_tmp9467 = 32'sh0000042e;
	assign w_sys_tmp9472 = (w_sys_tmp9473 + r_run_k_29);
	assign w_sys_tmp9473 = 32'sh00000493;
	assign w_sys_tmp9478 = (w_sys_tmp9479 + r_run_k_29);
	assign w_sys_tmp9479 = 32'sh000004f8;
	assign w_sys_tmp9484 = (w_sys_tmp9485 + r_run_k_29);
	assign w_sys_tmp9485 = 32'sh0000055d;
	assign w_sys_tmp9490 = (w_sys_tmp9491 + r_run_k_29);
	assign w_sys_tmp9491 = 32'sh000005c2;
	assign w_sys_tmp9496 = (w_sys_tmp9497 + r_run_k_29);
	assign w_sys_tmp9497 = 32'sh00000627;
	assign w_sys_tmp9502 = (w_sys_tmp9503 + r_run_k_29);
	assign w_sys_tmp9503 = 32'sh0000068c;
	assign w_sys_tmp9508 = (w_sys_tmp9509 + r_run_k_29);
	assign w_sys_tmp9509 = 32'sh000006f1;
	assign w_sys_tmp9514 = (w_sys_tmp9515 + r_run_k_29);
	assign w_sys_tmp9515 = 32'sh00000756;
	assign w_sys_tmp9520 = (w_sys_tmp9521 + r_run_k_29);
	assign w_sys_tmp9521 = 32'sh000007bb;
	assign w_sys_tmp9526 = (w_sys_tmp9527 + r_run_k_29);
	assign w_sys_tmp9527 = 32'sh00000820;
	assign w_sys_tmp9532 = (w_sys_tmp9533 + r_run_k_29);
	assign w_sys_tmp9533 = 32'sh00000885;
	assign w_sys_tmp9538 = (w_sys_tmp9539 + r_run_k_29);
	assign w_sys_tmp9539 = 32'sh000008ea;
	assign w_sys_tmp9556 = (w_sys_tmp9557 + r_run_k_29);
	assign w_sys_tmp9557 = 32'sh0000094f;
	assign w_sys_tmp9562 = (w_sys_tmp9563 + r_run_k_29);
	assign w_sys_tmp9563 = 32'sh000009b4;
	assign w_sys_tmp9568 = (w_sys_tmp9569 + r_run_k_29);
	assign w_sys_tmp9569 = 32'sh00000a19;
	assign w_sys_tmp9574 = (w_sys_tmp9575 + r_run_k_29);
	assign w_sys_tmp9575 = 32'sh00000a7e;
	assign w_sys_tmp9580 = (w_sys_tmp9581 + r_run_k_29);
	assign w_sys_tmp9581 = 32'sh00000ae3;
	assign w_sys_tmp9586 = (w_sys_tmp9587 + r_run_k_29);
	assign w_sys_tmp9587 = 32'sh00000b48;
	assign w_sys_tmp9592 = (w_sys_tmp9593 + r_run_k_29);
	assign w_sys_tmp9593 = 32'sh00000bad;
	assign w_sys_tmp9598 = (w_sys_tmp9599 + r_run_k_29);
	assign w_sys_tmp9599 = 32'sh00000c12;
	assign w_sys_tmp9604 = (w_sys_tmp9605 + r_run_k_29);
	assign w_sys_tmp9605 = 32'sh00000c77;
	assign w_sys_tmp9610 = (w_sys_tmp9611 + r_run_k_29);
	assign w_sys_tmp9611 = 32'sh00000cdc;
	assign w_sys_tmp9616 = (w_sys_tmp9617 + r_run_k_29);
	assign w_sys_tmp9617 = 32'sh00000d41;
	assign w_sys_tmp9622 = (w_sys_tmp9623 + r_run_k_29);
	assign w_sys_tmp9623 = 32'sh00000da6;
	assign w_sys_tmp9628 = (w_sys_tmp9629 + r_run_k_29);
	assign w_sys_tmp9629 = 32'sh00000e0b;
	assign w_sys_tmp9634 = (w_sys_tmp9635 + r_run_k_29);
	assign w_sys_tmp9635 = 32'sh00000e70;
	assign w_sys_tmp9640 = (w_sys_tmp9641 + r_run_k_29);
	assign w_sys_tmp9641 = 32'sh00000ed5;
	assign w_sys_tmp9646 = (w_sys_tmp9647 + r_run_k_29);
	assign w_sys_tmp9647 = 32'sh00000f3a;
	assign w_sys_tmp9652 = (w_sys_tmp9653 + r_run_k_29);
	assign w_sys_tmp9653 = 32'sh00000f9f;
	assign w_sys_tmp9658 = (w_sys_tmp9659 + r_run_k_29);
	assign w_sys_tmp9659 = 32'sh00001004;
	assign w_sys_tmp9664 = (w_sys_tmp9665 + r_run_k_29);
	assign w_sys_tmp9665 = 32'sh00001069;
	assign w_sys_tmp9670 = (w_sys_tmp9671 + r_run_k_29);
	assign w_sys_tmp9671 = 32'sh000010ce;
	assign w_sys_tmp9688 = (w_sys_tmp9689 + r_run_k_29);
	assign w_sys_tmp9689 = 32'sh00001133;
	assign w_sys_tmp9694 = (w_sys_tmp9695 + r_run_k_29);
	assign w_sys_tmp9695 = 32'sh00001198;
	assign w_sys_tmp9700 = (w_sys_tmp9701 + r_run_k_29);
	assign w_sys_tmp9701 = 32'sh000011fd;
	assign w_sys_tmp9706 = (w_sys_tmp9707 + r_run_k_29);
	assign w_sys_tmp9707 = 32'sh00001262;
	assign w_sys_tmp9712 = (w_sys_tmp9713 + r_run_k_29);
	assign w_sys_tmp9713 = 32'sh000012c7;
	assign w_sys_tmp9718 = (w_sys_tmp9719 + r_run_k_29);
	assign w_sys_tmp9719 = 32'sh000196ac;
	assign w_sys_tmp9724 = (w_sys_tmp9725 + r_run_k_29);
	assign w_sys_tmp9725 = 32'sh00001391;
	assign w_sys_tmp9730 = (w_sys_tmp9731 + r_run_k_29);
	assign w_sys_tmp9731 = 32'sh000013f6;
	assign w_sys_tmp9736 = (w_sys_tmp9737 + r_run_k_29);
	assign w_sys_tmp9737 = 32'sh0000145b;
	assign w_sys_tmp9742 = (w_sys_tmp9743 + r_run_k_29);
	assign w_sys_tmp9743 = 32'sh000014c0;
	assign w_sys_tmp9748 = (w_sys_tmp9749 + r_run_k_29);
	assign w_sys_tmp9749 = 32'sh00001525;
	assign w_sys_tmp9754 = (w_sys_tmp9755 + r_run_k_29);
	assign w_sys_tmp9755 = 32'sh0000158a;
	assign w_sys_tmp9760 = (w_sys_tmp9761 + r_run_k_29);
	assign w_sys_tmp9761 = 32'sh000015ef;
	assign w_sys_tmp9766 = (w_sys_tmp9767 + r_run_k_29);
	assign w_sys_tmp9767 = 32'sh00001654;
	assign w_sys_tmp9772 = (w_sys_tmp9773 + r_run_k_29);
	assign w_sys_tmp9773 = 32'sh000016b9;
	assign w_sys_tmp9778 = (w_sys_tmp9779 + r_run_k_29);
	assign w_sys_tmp9779 = 32'sh0000171e;
	assign w_sys_tmp9784 = (w_sys_tmp9785 + r_run_k_29);
	assign w_sys_tmp9785 = 32'sh00001783;
	assign w_sys_tmp9790 = (w_sys_tmp9791 + r_run_k_29);
	assign w_sys_tmp9791 = 32'sh000017e8;
	assign w_sys_tmp9796 = (w_sys_tmp9797 + r_run_k_29);
	assign w_sys_tmp9797 = 32'sh0000184d;
	assign w_sys_tmp9802 = (w_sys_tmp9803 + r_run_k_29);
	assign w_sys_tmp9803 = 32'sh000018b2;
	assign w_sys_tmp9820 = (w_sys_tmp9821 + r_run_k_29);
	assign w_sys_tmp9821 = 32'sh00001917;
	assign w_sys_tmp9826 = (w_sys_tmp9827 + r_run_k_29);
	assign w_sys_tmp9827 = 32'sh0000197c;
	assign w_sys_tmp9832 = (w_sys_tmp9833 + r_run_k_29);
	assign w_sys_tmp9833 = 32'sh000019e1;
	assign w_sys_tmp9838 = (w_sys_tmp9839 + r_run_k_29);
	assign w_sys_tmp9839 = 32'sh00001a46;
	assign w_sys_tmp9844 = (w_sys_tmp9845 + r_run_k_29);
	assign w_sys_tmp9845 = 32'sh00001aab;
	assign w_sys_tmp9850 = (w_sys_tmp9851 + r_run_k_29);
	assign w_sys_tmp9851 = 32'sh00001b10;
	assign w_sys_tmp9856 = (w_sys_tmp9857 + r_run_k_29);
	assign w_sys_tmp9857 = 32'sh00001b75;
	assign w_sys_tmp9862 = (w_sys_tmp9863 + r_run_k_29);
	assign w_sys_tmp9863 = 32'sh00001bda;
	assign w_sys_tmp9868 = (w_sys_tmp9869 + r_run_k_29);
	assign w_sys_tmp9869 = 32'sh00001c3f;
	assign w_sys_tmp9874 = (w_sys_tmp9875 + r_run_k_29);
	assign w_sys_tmp9875 = 32'sh00001ca4;
	assign w_sys_tmp9880 = (w_sys_tmp9881 + r_run_k_29);
	assign w_sys_tmp9881 = 32'sh00001d09;
	assign w_sys_tmp9886 = (w_sys_tmp9887 + r_run_k_29);
	assign w_sys_tmp9887 = 32'sh00001d6e;
	assign w_sys_tmp9892 = (w_sys_tmp9893 + r_run_k_29);
	assign w_sys_tmp9893 = 32'sh00001dd3;
	assign w_sys_tmp9898 = (w_sys_tmp9899 + r_run_k_29);
	assign w_sys_tmp9899 = 32'sh00001e38;
	assign w_sys_tmp9904 = (w_sys_tmp9905 + r_run_k_29);
	assign w_sys_tmp9905 = 32'sh00001e9d;
	assign w_sys_tmp9910 = (w_sys_tmp9911 + r_run_k_29);
	assign w_sys_tmp9911 = 32'sh00001f02;
	assign w_sys_tmp9916 = (w_sys_tmp9917 + r_run_k_29);
	assign w_sys_tmp9917 = 32'sh00001f67;
	assign w_sys_tmp9922 = (w_sys_tmp9923 + r_run_k_29);
	assign w_sys_tmp9923 = 32'sh00001fcc;
	assign w_sys_tmp9928 = (w_sys_tmp9929 + r_run_k_29);
	assign w_sys_tmp9929 = 32'sh00002031;
	assign w_sys_tmp9934 = (w_sys_tmp9935 + r_run_k_29);
	assign w_sys_tmp9935 = 32'sh00002096;
	assign w_sys_tmp9952 = (w_sys_tmp9953 + r_run_k_29);
	assign w_sys_tmp9953 = 32'sh000020fb;
	assign w_sys_tmp9958 = (w_sys_tmp9959 + r_run_k_29);
	assign w_sys_tmp9959 = 32'sh000c5de0;
	assign w_sys_tmp9964 = (w_sys_tmp9965 + r_run_k_29);
	assign w_sys_tmp9965 = 32'sh000021c5;
	assign w_sys_tmp9970 = (w_sys_tmp9971 + r_run_k_29);
	assign w_sys_tmp9971 = 32'sh0000222a;
	assign w_sys_tmp9976 = (w_sys_tmp9977 + r_run_k_29);
	assign w_sys_tmp9977 = 32'sh0000228f;
	assign w_sys_tmp9982 = (w_sys_tmp9983 + r_run_k_29);
	assign w_sys_tmp9983 = 32'sh000022f4;
	assign w_sys_tmp9988 = (w_sys_tmp9989 + r_run_k_29);
	assign w_sys_tmp9989 = 32'sh00002359;
	assign w_sys_tmp9994 = (w_sys_tmp9995 + r_run_k_29);
	assign w_sys_tmp9995 = 32'sh000023be;
	assign w_sys_tmp10000 = (w_sys_tmp10001 + r_run_k_29);
	assign w_sys_tmp10001 = 32'sh00002423;
	assign w_sys_tmp10006 = (w_sys_tmp10007 + r_run_k_29);
	assign w_sys_tmp10007 = 32'sh00002488;
	assign w_sys_tmp10012 = (w_sys_tmp10013 + r_run_k_29);
	assign w_sys_tmp10013 = 32'sh000024ed;
	assign w_sys_tmp10018 = (w_sys_tmp10019 + r_run_k_29);
	assign w_sys_tmp10019 = 32'sh00002552;
	assign w_sys_tmp10024 = (w_sys_tmp10025 + r_run_k_29);
	assign w_sys_tmp10025 = 32'sh000025b7;
	assign w_sys_tmp10030 = (w_sys_tmp10031 + r_run_k_29);
	assign w_sys_tmp10031 = 32'sh0000261c;
	assign w_sys_tmp10036 = (w_sys_tmp10037 + r_run_k_29);
	assign w_sys_tmp10037 = 32'sh00002681;
	assign w_sys_tmp10042 = (w_sys_tmp10043 + r_run_k_29);
	assign w_sys_tmp10043 = 32'sh000026e6;
	assign w_sys_tmp10048 = (w_sys_tmp10049 + r_run_k_29);
	assign w_sys_tmp10049 = 32'sh0000274b;
	assign w_sys_tmp10054 = (w_sys_tmp10055 + r_run_k_29);
	assign w_sys_tmp10055 = 32'sh000027b0;
	assign w_sys_tmp10060 = (w_sys_tmp10061 + r_run_k_29);
	assign w_sys_tmp10061 = 32'sh00002815;
	assign w_sys_tmp10065 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp10066 = 32'sh00000051;
	assign w_sys_tmp10067 = ( !w_sys_tmp10068 );
	assign w_sys_tmp10068 = (w_sys_tmp10069 < r_run_k_29);
	assign w_sys_tmp10069 = 32'sh00000065;
	assign w_sys_tmp10072 = (w_sys_tmp10073 + r_run_k_29);
	assign w_sys_tmp10073 = 32'sh00000065;
	assign w_sys_tmp10074 = w_fld_T_0_dataout_1;
	assign w_sys_tmp10078 = (w_sys_tmp10079 + r_run_k_29);
	assign w_sys_tmp10079 = 32'sh000000ca;
	assign w_sys_tmp10084 = (w_sys_tmp10085 + r_run_k_29);
	assign w_sys_tmp10085 = 32'sh0000012f;
	assign w_sys_tmp10090 = (w_sys_tmp10091 + r_run_k_29);
	assign w_sys_tmp10091 = 32'sh00000194;
	assign w_sys_tmp10096 = (w_sys_tmp10097 + r_run_k_29);
	assign w_sys_tmp10097 = 32'sh000001f9;
	assign w_sys_tmp10102 = (w_sys_tmp10103 + r_run_k_29);
	assign w_sys_tmp10103 = 32'sh0000025e;
	assign w_sys_tmp10108 = (w_sys_tmp10109 + r_run_k_29);
	assign w_sys_tmp10109 = 32'sh000002c3;
	assign w_sys_tmp10114 = (w_sys_tmp10115 + r_run_k_29);
	assign w_sys_tmp10115 = 32'sh00000328;
	assign w_sys_tmp10120 = (w_sys_tmp10121 + r_run_k_29);
	assign w_sys_tmp10121 = 32'sh0000038d;
	assign w_sys_tmp10126 = (w_sys_tmp10127 + r_run_k_29);
	assign w_sys_tmp10127 = 32'sh000003f2;
	assign w_sys_tmp10132 = (w_sys_tmp10133 + r_run_k_29);
	assign w_sys_tmp10133 = 32'sh00000457;
	assign w_sys_tmp10138 = (w_sys_tmp10139 + r_run_k_29);
	assign w_sys_tmp10139 = 32'sh000004bc;
	assign w_sys_tmp10144 = (w_sys_tmp10145 + r_run_k_29);
	assign w_sys_tmp10145 = 32'sh00000521;
	assign w_sys_tmp10150 = (w_sys_tmp10151 + r_run_k_29);
	assign w_sys_tmp10151 = 32'sh00000586;
	assign w_sys_tmp10156 = (w_sys_tmp10157 + r_run_k_29);
	assign w_sys_tmp10157 = 32'sh000005eb;
	assign w_sys_tmp10162 = (w_sys_tmp10163 + r_run_k_29);
	assign w_sys_tmp10163 = 32'sh00000650;
	assign w_sys_tmp10168 = (w_sys_tmp10169 + r_run_k_29);
	assign w_sys_tmp10169 = 32'sh000006b5;
	assign w_sys_tmp10174 = (w_sys_tmp10175 + r_run_k_29);
	assign w_sys_tmp10175 = 32'sh0000071a;
	assign w_sys_tmp10180 = (w_sys_tmp10181 + r_run_k_29);
	assign w_sys_tmp10181 = 32'sh0000077f;
	assign w_sys_tmp10186 = (w_sys_tmp10187 + r_run_k_29);
	assign w_sys_tmp10187 = 32'sh000007e4;
	assign w_sys_tmp10192 = (w_sys_tmp10193 + r_run_k_29);
	assign w_sys_tmp10193 = 32'sh00000849;
	assign w_sys_tmp10198 = (w_sys_tmp10199 + r_run_k_29);
	assign w_sys_tmp10199 = 32'sh000008ae;
	assign w_sys_tmp10216 = (w_sys_tmp10217 + r_run_k_29);
	assign w_sys_tmp10217 = 32'sh00000913;
	assign w_sys_tmp10222 = (w_sys_tmp10223 + r_run_k_29);
	assign w_sys_tmp10223 = 32'sh00000978;
	assign w_sys_tmp10228 = (w_sys_tmp10229 + r_run_k_29);
	assign w_sys_tmp10229 = 32'sh000009dd;
	assign w_sys_tmp10234 = (w_sys_tmp10235 + r_run_k_29);
	assign w_sys_tmp10235 = 32'sh00000a42;
	assign w_sys_tmp10240 = (w_sys_tmp10241 + r_run_k_29);
	assign w_sys_tmp10241 = 32'sh00000aa7;
	assign w_sys_tmp10246 = (w_sys_tmp10247 + r_run_k_29);
	assign w_sys_tmp10247 = 32'sh00000b0c;
	assign w_sys_tmp10252 = (w_sys_tmp10253 + r_run_k_29);
	assign w_sys_tmp10253 = 32'sh00000b71;
	assign w_sys_tmp10258 = (w_sys_tmp10259 + r_run_k_29);
	assign w_sys_tmp10259 = 32'sh00000bd6;
	assign w_sys_tmp10264 = (w_sys_tmp10265 + r_run_k_29);
	assign w_sys_tmp10265 = 32'sh00000c3b;
	assign w_sys_tmp10270 = (w_sys_tmp10271 + r_run_k_29);
	assign w_sys_tmp10271 = 32'sh00000ca0;
	assign w_sys_tmp10276 = (w_sys_tmp10277 + r_run_k_29);
	assign w_sys_tmp10277 = 32'sh00000d05;
	assign w_sys_tmp10282 = (w_sys_tmp10283 + r_run_k_29);
	assign w_sys_tmp10283 = 32'sh00000d6a;
	assign w_sys_tmp10288 = (w_sys_tmp10289 + r_run_k_29);
	assign w_sys_tmp10289 = 32'sh00000dcf;
	assign w_sys_tmp10294 = (w_sys_tmp10295 + r_run_k_29);
	assign w_sys_tmp10295 = 32'sh00000e34;
	assign w_sys_tmp10300 = (w_sys_tmp10301 + r_run_k_29);
	assign w_sys_tmp10301 = 32'sh00000e99;
	assign w_sys_tmp10306 = (w_sys_tmp10307 + r_run_k_29);
	assign w_sys_tmp10307 = 32'sh00000efe;
	assign w_sys_tmp10312 = (w_sys_tmp10313 + r_run_k_29);
	assign w_sys_tmp10313 = 32'sh00000f63;
	assign w_sys_tmp10318 = (w_sys_tmp10319 + r_run_k_29);
	assign w_sys_tmp10319 = 32'sh00000fc8;
	assign w_sys_tmp10324 = (w_sys_tmp10325 + r_run_k_29);
	assign w_sys_tmp10325 = 32'sh0000102d;
	assign w_sys_tmp10330 = (w_sys_tmp10331 + r_run_k_29);
	assign w_sys_tmp10331 = 32'sh00001092;
	assign w_sys_tmp10348 = (w_sys_tmp10349 + r_run_k_29);
	assign w_sys_tmp10349 = 32'sh000010f7;
	assign w_sys_tmp10354 = (w_sys_tmp10355 + r_run_k_29);
	assign w_sys_tmp10355 = 32'sh0000115c;
	assign w_sys_tmp10360 = (w_sys_tmp10361 + r_run_k_29);
	assign w_sys_tmp10361 = 32'sh000011c1;
	assign w_sys_tmp10366 = (w_sys_tmp10367 + r_run_k_29);
	assign w_sys_tmp10367 = 32'sh00001226;
	assign w_sys_tmp10372 = (w_sys_tmp10373 + r_run_k_29);
	assign w_sys_tmp10373 = 32'sh0000128b;
	assign w_sys_tmp10378 = (w_sys_tmp10379 + r_run_k_29);
	assign w_sys_tmp10379 = 32'sh00019670;
	assign w_sys_tmp10384 = (w_sys_tmp10385 + r_run_k_29);
	assign w_sys_tmp10385 = 32'sh00001355;
	assign w_sys_tmp10390 = (w_sys_tmp10391 + r_run_k_29);
	assign w_sys_tmp10391 = 32'sh000013ba;
	assign w_sys_tmp10396 = (w_sys_tmp10397 + r_run_k_29);
	assign w_sys_tmp10397 = 32'sh0000141f;
	assign w_sys_tmp10402 = (w_sys_tmp10403 + r_run_k_29);
	assign w_sys_tmp10403 = 32'sh00001484;
	assign w_sys_tmp10408 = (w_sys_tmp10409 + r_run_k_29);
	assign w_sys_tmp10409 = 32'sh000014e9;
	assign w_sys_tmp10414 = (w_sys_tmp10415 + r_run_k_29);
	assign w_sys_tmp10415 = 32'sh0000154e;
	assign w_sys_tmp10420 = (w_sys_tmp10421 + r_run_k_29);
	assign w_sys_tmp10421 = 32'sh000015b3;
	assign w_sys_tmp10426 = (w_sys_tmp10427 + r_run_k_29);
	assign w_sys_tmp10427 = 32'sh00001618;
	assign w_sys_tmp10432 = (w_sys_tmp10433 + r_run_k_29);
	assign w_sys_tmp10433 = 32'sh0000167d;
	assign w_sys_tmp10438 = (w_sys_tmp10439 + r_run_k_29);
	assign w_sys_tmp10439 = 32'sh000016e2;
	assign w_sys_tmp10444 = (w_sys_tmp10445 + r_run_k_29);
	assign w_sys_tmp10445 = 32'sh00001747;
	assign w_sys_tmp10450 = (w_sys_tmp10451 + r_run_k_29);
	assign w_sys_tmp10451 = 32'sh000017ac;
	assign w_sys_tmp10456 = (w_sys_tmp10457 + r_run_k_29);
	assign w_sys_tmp10457 = 32'sh00001811;
	assign w_sys_tmp10462 = (w_sys_tmp10463 + r_run_k_29);
	assign w_sys_tmp10463 = 32'sh00001876;
	assign w_sys_tmp10480 = (w_sys_tmp10481 + r_run_k_29);
	assign w_sys_tmp10481 = 32'sh000018db;
	assign w_sys_tmp10486 = (w_sys_tmp10487 + r_run_k_29);
	assign w_sys_tmp10487 = 32'sh00001940;
	assign w_sys_tmp10492 = (w_sys_tmp10493 + r_run_k_29);
	assign w_sys_tmp10493 = 32'sh000019a5;
	assign w_sys_tmp10498 = (w_sys_tmp10499 + r_run_k_29);
	assign w_sys_tmp10499 = 32'sh00001a0a;
	assign w_sys_tmp10504 = (w_sys_tmp10505 + r_run_k_29);
	assign w_sys_tmp10505 = 32'sh00001a6f;
	assign w_sys_tmp10510 = (w_sys_tmp10511 + r_run_k_29);
	assign w_sys_tmp10511 = 32'sh00001ad4;
	assign w_sys_tmp10516 = (w_sys_tmp10517 + r_run_k_29);
	assign w_sys_tmp10517 = 32'sh00001b39;
	assign w_sys_tmp10522 = (w_sys_tmp10523 + r_run_k_29);
	assign w_sys_tmp10523 = 32'sh00001b9e;
	assign w_sys_tmp10528 = (w_sys_tmp10529 + r_run_k_29);
	assign w_sys_tmp10529 = 32'sh00001c03;
	assign w_sys_tmp10534 = (w_sys_tmp10535 + r_run_k_29);
	assign w_sys_tmp10535 = 32'sh00001c68;
	assign w_sys_tmp10540 = (w_sys_tmp10541 + r_run_k_29);
	assign w_sys_tmp10541 = 32'sh00001ccd;
	assign w_sys_tmp10546 = (w_sys_tmp10547 + r_run_k_29);
	assign w_sys_tmp10547 = 32'sh00001d32;
	assign w_sys_tmp10552 = (w_sys_tmp10553 + r_run_k_29);
	assign w_sys_tmp10553 = 32'sh00001d97;
	assign w_sys_tmp10558 = (w_sys_tmp10559 + r_run_k_29);
	assign w_sys_tmp10559 = 32'sh00001dfc;
	assign w_sys_tmp10564 = (w_sys_tmp10565 + r_run_k_29);
	assign w_sys_tmp10565 = 32'sh00001e61;
	assign w_sys_tmp10570 = (w_sys_tmp10571 + r_run_k_29);
	assign w_sys_tmp10571 = 32'sh00001ec6;
	assign w_sys_tmp10576 = (w_sys_tmp10577 + r_run_k_29);
	assign w_sys_tmp10577 = 32'sh00001f2b;
	assign w_sys_tmp10582 = (w_sys_tmp10583 + r_run_k_29);
	assign w_sys_tmp10583 = 32'sh00001f90;
	assign w_sys_tmp10588 = (w_sys_tmp10589 + r_run_k_29);
	assign w_sys_tmp10589 = 32'sh00001ff5;
	assign w_sys_tmp10594 = (w_sys_tmp10595 + r_run_k_29);
	assign w_sys_tmp10595 = 32'sh0000205a;
	assign w_sys_tmp10612 = (w_sys_tmp10613 + r_run_k_29);
	assign w_sys_tmp10613 = 32'sh000020bf;
	assign w_sys_tmp10618 = (w_sys_tmp10619 + r_run_k_29);
	assign w_sys_tmp10619 = 32'sh000c5da4;
	assign w_sys_tmp10624 = (w_sys_tmp10625 + r_run_k_29);
	assign w_sys_tmp10625 = 32'sh00002189;
	assign w_sys_tmp10630 = (w_sys_tmp10631 + r_run_k_29);
	assign w_sys_tmp10631 = 32'sh000021ee;
	assign w_sys_tmp10636 = (w_sys_tmp10637 + r_run_k_29);
	assign w_sys_tmp10637 = 32'sh00002253;
	assign w_sys_tmp10642 = (w_sys_tmp10643 + r_run_k_29);
	assign w_sys_tmp10643 = 32'sh000022b8;
	assign w_sys_tmp10648 = (w_sys_tmp10649 + r_run_k_29);
	assign w_sys_tmp10649 = 32'sh0000231d;
	assign w_sys_tmp10654 = (w_sys_tmp10655 + r_run_k_29);
	assign w_sys_tmp10655 = 32'sh00002382;
	assign w_sys_tmp10660 = (w_sys_tmp10661 + r_run_k_29);
	assign w_sys_tmp10661 = 32'sh000023e7;
	assign w_sys_tmp10666 = (w_sys_tmp10667 + r_run_k_29);
	assign w_sys_tmp10667 = 32'sh0000244c;
	assign w_sys_tmp10672 = (w_sys_tmp10673 + r_run_k_29);
	assign w_sys_tmp10673 = 32'sh000024b1;
	assign w_sys_tmp10678 = (w_sys_tmp10679 + r_run_k_29);
	assign w_sys_tmp10679 = 32'sh00002516;
	assign w_sys_tmp10684 = (w_sys_tmp10685 + r_run_k_29);
	assign w_sys_tmp10685 = 32'sh0000257b;
	assign w_sys_tmp10690 = (w_sys_tmp10691 + r_run_k_29);
	assign w_sys_tmp10691 = 32'sh000025e0;
	assign w_sys_tmp10696 = (w_sys_tmp10697 + r_run_k_29);
	assign w_sys_tmp10697 = 32'sh00002645;
	assign w_sys_tmp10702 = (w_sys_tmp10703 + r_run_k_29);
	assign w_sys_tmp10703 = 32'sh000026aa;
	assign w_sys_tmp10708 = (w_sys_tmp10709 + r_run_k_29);
	assign w_sys_tmp10709 = 32'sh0000270f;
	assign w_sys_tmp10714 = (w_sys_tmp10715 + r_run_k_29);
	assign w_sys_tmp10715 = 32'sh00002774;
	assign w_sys_tmp10720 = (w_sys_tmp10721 + r_run_k_29);
	assign w_sys_tmp10721 = 32'sh000027d9;
	assign w_sys_tmp10725 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp10726 = 32'sh00000002;
	assign w_sys_tmp10727 = ( !w_sys_tmp10728 );
	assign w_sys_tmp10728 = (w_sys_tmp10729 < r_run_k_29);
	assign w_sys_tmp10729 = 32'sh00000015;
	assign w_sys_tmp10732 = (w_sys_tmp10733 + r_run_k_29);
	assign w_sys_tmp10733 = 32'sh000000ca;
	assign w_sys_tmp10734 = w_sub00_result_dataout;
	assign w_sys_tmp10738 = (w_sys_tmp10739 + r_run_k_29);
	assign w_sys_tmp10739 = 32'sh0000012f;
	assign w_sys_tmp10744 = (w_sys_tmp10745 + r_run_k_29);
	assign w_sys_tmp10745 = 32'sh00000194;
	assign w_sys_tmp10750 = (w_sys_tmp10751 + r_run_k_29);
	assign w_sys_tmp10751 = 32'sh000001f9;
	assign w_sys_tmp10756 = (w_sys_tmp10757 + r_run_k_29);
	assign w_sys_tmp10757 = 32'sh0000025e;
	assign w_sys_tmp10762 = (w_sys_tmp10763 + r_run_k_29);
	assign w_sys_tmp10763 = 32'sh000002c3;
	assign w_sys_tmp10768 = (w_sys_tmp10769 + r_run_k_29);
	assign w_sys_tmp10769 = 32'sh00000328;
	assign w_sys_tmp10774 = (w_sys_tmp10775 + r_run_k_29);
	assign w_sys_tmp10775 = 32'sh0000038d;
	assign w_sys_tmp10780 = (w_sys_tmp10781 + r_run_k_29);
	assign w_sys_tmp10781 = 32'sh000003f2;
	assign w_sys_tmp10786 = (w_sys_tmp10787 + r_run_k_29);
	assign w_sys_tmp10787 = 32'sh00000457;
	assign w_sys_tmp10792 = (w_sys_tmp10793 + r_run_k_29);
	assign w_sys_tmp10793 = 32'sh000004bc;
	assign w_sys_tmp10798 = (w_sys_tmp10799 + r_run_k_29);
	assign w_sys_tmp10799 = 32'sh00000521;
	assign w_sys_tmp10804 = (w_sys_tmp10805 + r_run_k_29);
	assign w_sys_tmp10805 = 32'sh00000586;
	assign w_sys_tmp10810 = (w_sys_tmp10811 + r_run_k_29);
	assign w_sys_tmp10811 = 32'sh000005eb;
	assign w_sys_tmp10816 = (w_sys_tmp10817 + r_run_k_29);
	assign w_sys_tmp10817 = 32'sh00000650;
	assign w_sys_tmp10822 = (w_sys_tmp10823 + r_run_k_29);
	assign w_sys_tmp10823 = 32'sh000006b5;
	assign w_sys_tmp10828 = (w_sys_tmp10829 + r_run_k_29);
	assign w_sys_tmp10829 = 32'sh0000071a;
	assign w_sys_tmp10834 = (w_sys_tmp10835 + r_run_k_29);
	assign w_sys_tmp10835 = 32'sh0000077f;
	assign w_sys_tmp10840 = (w_sys_tmp10841 + r_run_k_29);
	assign w_sys_tmp10841 = 32'sh000007e4;
	assign w_sys_tmp10846 = (w_sys_tmp10847 + r_run_k_29);
	assign w_sys_tmp10847 = 32'sh00000849;
	assign w_sys_tmp10922 = (w_sys_tmp10923 + r_run_k_29);
	assign w_sys_tmp10923 = 32'sh000008ae;
	assign w_sys_tmp10927 = (w_sys_tmp10928 + r_run_k_29);
	assign w_sys_tmp10928 = 32'sh00000913;
	assign w_sys_tmp10932 = (w_sys_tmp10933 + r_run_k_29);
	assign w_sys_tmp10933 = 32'sh00000978;
	assign w_sys_tmp10937 = (w_sys_tmp10938 + r_run_k_29);
	assign w_sys_tmp10938 = 32'sh000009dd;
	assign w_sys_tmp10942 = (w_sys_tmp10943 + r_run_k_29);
	assign w_sys_tmp10943 = 32'sh00000a42;
	assign w_sys_tmp10947 = (w_sys_tmp10948 + r_run_k_29);
	assign w_sys_tmp10948 = 32'sh00000aa7;
	assign w_sys_tmp10952 = (w_sys_tmp10953 + r_run_k_29);
	assign w_sys_tmp10953 = 32'sh00000b0c;
	assign w_sys_tmp10957 = (w_sys_tmp10958 + r_run_k_29);
	assign w_sys_tmp10958 = 32'sh00000b71;
	assign w_sys_tmp10962 = (w_sys_tmp10963 + r_run_k_29);
	assign w_sys_tmp10963 = 32'sh00000bd6;
	assign w_sys_tmp10967 = (w_sys_tmp10968 + r_run_k_29);
	assign w_sys_tmp10968 = 32'sh00000c3b;
	assign w_sys_tmp10972 = (w_sys_tmp10973 + r_run_k_29);
	assign w_sys_tmp10973 = 32'sh00000ca0;
	assign w_sys_tmp10977 = (w_sys_tmp10978 + r_run_k_29);
	assign w_sys_tmp10978 = 32'sh00000d05;
	assign w_sys_tmp10982 = (w_sys_tmp10983 + r_run_k_29);
	assign w_sys_tmp10983 = 32'sh00000d6a;
	assign w_sys_tmp10987 = (w_sys_tmp10988 + r_run_k_29);
	assign w_sys_tmp10988 = 32'sh00000dcf;
	assign w_sys_tmp10992 = (w_sys_tmp10993 + r_run_k_29);
	assign w_sys_tmp10993 = 32'sh00000e34;
	assign w_sys_tmp10997 = (w_sys_tmp10998 + r_run_k_29);
	assign w_sys_tmp10998 = 32'sh00000e99;
	assign w_sys_tmp11002 = (w_sys_tmp11003 + r_run_k_29);
	assign w_sys_tmp11003 = 32'sh00000efe;
	assign w_sys_tmp11007 = (w_sys_tmp11008 + r_run_k_29);
	assign w_sys_tmp11008 = 32'sh00000f63;
	assign w_sys_tmp11012 = (w_sys_tmp11013 + r_run_k_29);
	assign w_sys_tmp11013 = 32'sh00000fc8;
	assign w_sys_tmp11017 = (w_sys_tmp11018 + r_run_k_29);
	assign w_sys_tmp11018 = 32'sh0000102d;
	assign w_sys_tmp11162 = (w_sys_tmp11163 + r_run_k_29);
	assign w_sys_tmp11163 = 32'sh00001092;
	assign w_sys_tmp11167 = (w_sys_tmp11168 + r_run_k_29);
	assign w_sys_tmp11168 = 32'sh000010f7;
	assign w_sys_tmp11172 = (w_sys_tmp11173 + r_run_k_29);
	assign w_sys_tmp11173 = 32'sh0000115c;
	assign w_sys_tmp11177 = (w_sys_tmp11178 + r_run_k_29);
	assign w_sys_tmp11178 = 32'sh000011c1;
	assign w_sys_tmp11182 = (w_sys_tmp11183 + r_run_k_29);
	assign w_sys_tmp11183 = 32'sh00001226;
	assign w_sys_tmp11187 = (w_sys_tmp11188 + r_run_k_29);
	assign w_sys_tmp11188 = 32'sh0000128b;
	assign w_sys_tmp11192 = (w_sys_tmp11193 + r_run_k_29);
	assign w_sys_tmp11193 = 32'sh000012f0;
	assign w_sys_tmp11197 = (w_sys_tmp11198 + r_run_k_29);
	assign w_sys_tmp11198 = 32'sh00001355;
	assign w_sys_tmp11202 = (w_sys_tmp11203 + r_run_k_29);
	assign w_sys_tmp11203 = 32'sh000013ba;
	assign w_sys_tmp11207 = (w_sys_tmp11208 + r_run_k_29);
	assign w_sys_tmp11208 = 32'sh0000141f;
	assign w_sys_tmp11212 = (w_sys_tmp11213 + r_run_k_29);
	assign w_sys_tmp11213 = 32'sh00001484;
	assign w_sys_tmp11217 = (w_sys_tmp11218 + r_run_k_29);
	assign w_sys_tmp11218 = 32'sh000014e9;
	assign w_sys_tmp11222 = (w_sys_tmp11223 + r_run_k_29);
	assign w_sys_tmp11223 = 32'sh0000154e;
	assign w_sys_tmp11227 = (w_sys_tmp11228 + r_run_k_29);
	assign w_sys_tmp11228 = 32'sh000015b3;
	assign w_sys_tmp11232 = (w_sys_tmp11233 + r_run_k_29);
	assign w_sys_tmp11233 = 32'sh00001618;
	assign w_sys_tmp11237 = (w_sys_tmp11238 + r_run_k_29);
	assign w_sys_tmp11238 = 32'sh0000167d;
	assign w_sys_tmp11242 = (w_sys_tmp11243 + r_run_k_29);
	assign w_sys_tmp11243 = 32'sh000016e2;
	assign w_sys_tmp11247 = (w_sys_tmp11248 + r_run_k_29);
	assign w_sys_tmp11248 = 32'sh00001747;
	assign w_sys_tmp11252 = (w_sys_tmp11253 + r_run_k_29);
	assign w_sys_tmp11253 = 32'sh000017ac;
	assign w_sys_tmp11257 = (w_sys_tmp11258 + r_run_k_29);
	assign w_sys_tmp11258 = 32'sh00001811;
	assign w_sys_tmp11267 = (w_sys_tmp11268 + r_run_k_29);
	assign w_sys_tmp11268 = 32'sh00001876;
	assign w_sys_tmp11272 = (w_sys_tmp11273 + r_run_k_29);
	assign w_sys_tmp11273 = 32'sh000018db;
	assign w_sys_tmp11277 = (w_sys_tmp11278 + r_run_k_29);
	assign w_sys_tmp11278 = 32'sh00001940;
	assign w_sys_tmp11282 = (w_sys_tmp11283 + r_run_k_29);
	assign w_sys_tmp11283 = 32'sh000019a5;
	assign w_sys_tmp11287 = (w_sys_tmp11288 + r_run_k_29);
	assign w_sys_tmp11288 = 32'sh00001a0a;
	assign w_sys_tmp11292 = (w_sys_tmp11293 + r_run_k_29);
	assign w_sys_tmp11293 = 32'sh00001a6f;
	assign w_sys_tmp11297 = (w_sys_tmp11298 + r_run_k_29);
	assign w_sys_tmp11298 = 32'sh00001ad4;
	assign w_sys_tmp11302 = (w_sys_tmp11303 + r_run_k_29);
	assign w_sys_tmp11303 = 32'sh00001b39;
	assign w_sys_tmp11307 = (w_sys_tmp11308 + r_run_k_29);
	assign w_sys_tmp11308 = 32'sh00001b9e;
	assign w_sys_tmp11312 = (w_sys_tmp11313 + r_run_k_29);
	assign w_sys_tmp11313 = 32'sh00001c03;
	assign w_sys_tmp11317 = (w_sys_tmp11318 + r_run_k_29);
	assign w_sys_tmp11318 = 32'sh00001c68;
	assign w_sys_tmp11322 = (w_sys_tmp11323 + r_run_k_29);
	assign w_sys_tmp11323 = 32'sh00001ccd;
	assign w_sys_tmp11327 = (w_sys_tmp11328 + r_run_k_29);
	assign w_sys_tmp11328 = 32'sh00001d32;
	assign w_sys_tmp11332 = (w_sys_tmp11333 + r_run_k_29);
	assign w_sys_tmp11333 = 32'sh00001d97;
	assign w_sys_tmp11337 = (w_sys_tmp11338 + r_run_k_29);
	assign w_sys_tmp11338 = 32'sh00001dfc;
	assign w_sys_tmp11342 = (w_sys_tmp11343 + r_run_k_29);
	assign w_sys_tmp11343 = 32'sh00001e61;
	assign w_sys_tmp11347 = (w_sys_tmp11348 + r_run_k_29);
	assign w_sys_tmp11348 = 32'sh00001ec6;
	assign w_sys_tmp11352 = (w_sys_tmp11353 + r_run_k_29);
	assign w_sys_tmp11353 = 32'sh00001f2b;
	assign w_sys_tmp11357 = (w_sys_tmp11358 + r_run_k_29);
	assign w_sys_tmp11358 = 32'sh00001f90;
	assign w_sys_tmp11362 = (w_sys_tmp11363 + r_run_k_29);
	assign w_sys_tmp11363 = 32'sh00001ff5;
	assign w_sys_tmp11372 = (w_sys_tmp11373 + r_run_k_29);
	assign w_sys_tmp11373 = 32'sh0000205a;
	assign w_sys_tmp11377 = (w_sys_tmp11378 + r_run_k_29);
	assign w_sys_tmp11378 = 32'sh000020bf;
	assign w_sys_tmp11382 = (w_sys_tmp11383 + r_run_k_29);
	assign w_sys_tmp11383 = 32'sh00002124;
	assign w_sys_tmp11387 = (w_sys_tmp11388 + r_run_k_29);
	assign w_sys_tmp11388 = 32'sh00002189;
	assign w_sys_tmp11392 = (w_sys_tmp11393 + r_run_k_29);
	assign w_sys_tmp11393 = 32'sh000021ee;
	assign w_sys_tmp11397 = (w_sys_tmp11398 + r_run_k_29);
	assign w_sys_tmp11398 = 32'sh00002253;
	assign w_sys_tmp11402 = (w_sys_tmp11403 + r_run_k_29);
	assign w_sys_tmp11403 = 32'sh000022b8;
	assign w_sys_tmp11407 = (w_sys_tmp11408 + r_run_k_29);
	assign w_sys_tmp11408 = 32'sh0000231d;
	assign w_sys_tmp11412 = (w_sys_tmp11413 + r_run_k_29);
	assign w_sys_tmp11413 = 32'sh00002382;
	assign w_sys_tmp11417 = (w_sys_tmp11418 + r_run_k_29);
	assign w_sys_tmp11418 = 32'sh000023e7;
	assign w_sys_tmp11422 = (w_sys_tmp11423 + r_run_k_29);
	assign w_sys_tmp11423 = 32'sh0000244c;
	assign w_sys_tmp11427 = (w_sys_tmp11428 + r_run_k_29);
	assign w_sys_tmp11428 = 32'sh000024b1;
	assign w_sys_tmp11432 = (w_sys_tmp11433 + r_run_k_29);
	assign w_sys_tmp11433 = 32'sh00002516;
	assign w_sys_tmp11437 = (w_sys_tmp11438 + r_run_k_29);
	assign w_sys_tmp11438 = 32'sh0000257b;
	assign w_sys_tmp11442 = (w_sys_tmp11443 + r_run_k_29);
	assign w_sys_tmp11443 = 32'sh000025e0;
	assign w_sys_tmp11447 = (w_sys_tmp11448 + r_run_k_29);
	assign w_sys_tmp11448 = 32'sh00002645;
	assign w_sys_tmp11452 = (w_sys_tmp11453 + r_run_k_29);
	assign w_sys_tmp11453 = 32'sh000026aa;
	assign w_sys_tmp11457 = (w_sys_tmp11458 + r_run_k_29);
	assign w_sys_tmp11458 = 32'sh0000270f;
	assign w_sys_tmp11462 = (w_sys_tmp11463 + r_run_k_29);
	assign w_sys_tmp11463 = 32'sh00002774;
	assign w_sys_tmp11467 = (w_sys_tmp11468 + r_run_k_29);
	assign w_sys_tmp11468 = 32'sh000000de;
	assign w_sys_tmp11472 = (w_sys_tmp11473 + r_run_k_29);
	assign w_sys_tmp11473 = 32'sh00000143;
	assign w_sys_tmp11477 = (w_sys_tmp11478 + r_run_k_29);
	assign w_sys_tmp11478 = 32'sh000001a8;
	assign w_sys_tmp11482 = (w_sys_tmp11483 + r_run_k_29);
	assign w_sys_tmp11483 = 32'sh0000020d;
	assign w_sys_tmp11487 = (w_sys_tmp11488 + r_run_k_29);
	assign w_sys_tmp11488 = 32'sh00000272;
	assign w_sys_tmp11492 = (w_sys_tmp11493 + r_run_k_29);
	assign w_sys_tmp11493 = 32'sh000002d7;
	assign w_sys_tmp11497 = (w_sys_tmp11498 + r_run_k_29);
	assign w_sys_tmp11498 = 32'sh0000033c;
	assign w_sys_tmp11502 = (w_sys_tmp11503 + r_run_k_29);
	assign w_sys_tmp11503 = 32'sh000003a1;
	assign w_sys_tmp11507 = (w_sys_tmp11508 + r_run_k_29);
	assign w_sys_tmp11508 = 32'sh00000406;
	assign w_sys_tmp11512 = (w_sys_tmp11513 + r_run_k_29);
	assign w_sys_tmp11513 = 32'sh0000046b;
	assign w_sys_tmp11517 = (w_sys_tmp11518 + r_run_k_29);
	assign w_sys_tmp11518 = 32'sh000004d0;
	assign w_sys_tmp11522 = (w_sys_tmp11523 + r_run_k_29);
	assign w_sys_tmp11523 = 32'sh00000535;
	assign w_sys_tmp11527 = (w_sys_tmp11528 + r_run_k_29);
	assign w_sys_tmp11528 = 32'sh0000059a;
	assign w_sys_tmp11532 = (w_sys_tmp11533 + r_run_k_29);
	assign w_sys_tmp11533 = 32'sh000005ff;
	assign w_sys_tmp11537 = (w_sys_tmp11538 + r_run_k_29);
	assign w_sys_tmp11538 = 32'sh00000664;
	assign w_sys_tmp11542 = (w_sys_tmp11543 + r_run_k_29);
	assign w_sys_tmp11543 = 32'sh000006c9;
	assign w_sys_tmp11547 = (w_sys_tmp11548 + r_run_k_29);
	assign w_sys_tmp11548 = 32'sh0000072e;
	assign w_sys_tmp11552 = (w_sys_tmp11553 + r_run_k_29);
	assign w_sys_tmp11553 = 32'sh00000793;
	assign w_sys_tmp11557 = (w_sys_tmp11558 + r_run_k_29);
	assign w_sys_tmp11558 = 32'sh000007f8;
	assign w_sys_tmp11562 = (w_sys_tmp11563 + r_run_k_29);
	assign w_sys_tmp11563 = 32'sh0000085d;
	assign w_sys_tmp11567 = (w_sys_tmp11568 + r_run_k_29);
	assign w_sys_tmp11568 = 32'sh000008c2;
	assign w_sys_tmp11572 = (w_sys_tmp11573 + r_run_k_29);
	assign w_sys_tmp11573 = 32'sh00000927;
	assign w_sys_tmp11577 = (w_sys_tmp11578 + r_run_k_29);
	assign w_sys_tmp11578 = 32'sh0000098c;
	assign w_sys_tmp11582 = (w_sys_tmp11583 + r_run_k_29);
	assign w_sys_tmp11583 = 32'sh000009f1;
	assign w_sys_tmp11587 = (w_sys_tmp11588 + r_run_k_29);
	assign w_sys_tmp11588 = 32'sh00000a56;
	assign w_sys_tmp11592 = (w_sys_tmp11593 + r_run_k_29);
	assign w_sys_tmp11593 = 32'sh00000abb;
	assign w_sys_tmp11597 = (w_sys_tmp11598 + r_run_k_29);
	assign w_sys_tmp11598 = 32'sh00000b20;
	assign w_sys_tmp11602 = (w_sys_tmp11603 + r_run_k_29);
	assign w_sys_tmp11603 = 32'sh00000b85;
	assign w_sys_tmp11607 = (w_sys_tmp11608 + r_run_k_29);
	assign w_sys_tmp11608 = 32'sh00000bea;
	assign w_sys_tmp11612 = (w_sys_tmp11613 + r_run_k_29);
	assign w_sys_tmp11613 = 32'sh00000c4f;
	assign w_sys_tmp11617 = (w_sys_tmp11618 + r_run_k_29);
	assign w_sys_tmp11618 = 32'sh00000cb4;
	assign w_sys_tmp11622 = (w_sys_tmp11623 + r_run_k_29);
	assign w_sys_tmp11623 = 32'sh00000d19;
	assign w_sys_tmp11627 = (w_sys_tmp11628 + r_run_k_29);
	assign w_sys_tmp11628 = 32'sh00000d7e;
	assign w_sys_tmp11632 = (w_sys_tmp11633 + r_run_k_29);
	assign w_sys_tmp11633 = 32'sh00000de3;
	assign w_sys_tmp11637 = (w_sys_tmp11638 + r_run_k_29);
	assign w_sys_tmp11638 = 32'sh00000e48;
	assign w_sys_tmp11642 = (w_sys_tmp11643 + r_run_k_29);
	assign w_sys_tmp11643 = 32'sh00000ead;
	assign w_sys_tmp11647 = (w_sys_tmp11648 + r_run_k_29);
	assign w_sys_tmp11648 = 32'sh00000f12;
	assign w_sys_tmp11652 = (w_sys_tmp11653 + r_run_k_29);
	assign w_sys_tmp11653 = 32'sh00000f77;
	assign w_sys_tmp11657 = (w_sys_tmp11658 + r_run_k_29);
	assign w_sys_tmp11658 = 32'sh00000fdc;
	assign w_sys_tmp11662 = (w_sys_tmp11663 + r_run_k_29);
	assign w_sys_tmp11663 = 32'sh00001041;
	assign w_sys_tmp11667 = (w_sys_tmp11668 + r_run_k_29);
	assign w_sys_tmp11668 = 32'sh000010a6;
	assign w_sys_tmp11672 = (w_sys_tmp11673 + r_run_k_29);
	assign w_sys_tmp11673 = 32'sh0000110b;
	assign w_sys_tmp11677 = (w_sys_tmp11678 + r_run_k_29);
	assign w_sys_tmp11678 = 32'sh00001170;
	assign w_sys_tmp11682 = (w_sys_tmp11683 + r_run_k_29);
	assign w_sys_tmp11683 = 32'sh000011d5;
	assign w_sys_tmp11687 = (w_sys_tmp11688 + r_run_k_29);
	assign w_sys_tmp11688 = 32'sh0000123a;
	assign w_sys_tmp11692 = (w_sys_tmp11693 + r_run_k_29);
	assign w_sys_tmp11693 = 32'sh0000129f;
	assign w_sys_tmp11697 = (w_sys_tmp11698 + r_run_k_29);
	assign w_sys_tmp11698 = 32'sh00001304;
	assign w_sys_tmp11702 = (w_sys_tmp11703 + r_run_k_29);
	assign w_sys_tmp11703 = 32'sh00001369;
	assign w_sys_tmp11707 = (w_sys_tmp11708 + r_run_k_29);
	assign w_sys_tmp11708 = 32'sh000013ce;
	assign w_sys_tmp11712 = (w_sys_tmp11713 + r_run_k_29);
	assign w_sys_tmp11713 = 32'sh00001433;
	assign w_sys_tmp11717 = (w_sys_tmp11718 + r_run_k_29);
	assign w_sys_tmp11718 = 32'sh00001498;
	assign w_sys_tmp11722 = (w_sys_tmp11723 + r_run_k_29);
	assign w_sys_tmp11723 = 32'sh000014fd;
	assign w_sys_tmp11727 = (w_sys_tmp11728 + r_run_k_29);
	assign w_sys_tmp11728 = 32'sh00001562;
	assign w_sys_tmp11732 = (w_sys_tmp11733 + r_run_k_29);
	assign w_sys_tmp11733 = 32'sh000015c7;
	assign w_sys_tmp11737 = (w_sys_tmp11738 + r_run_k_29);
	assign w_sys_tmp11738 = 32'sh0000162c;
	assign w_sys_tmp11742 = (w_sys_tmp11743 + r_run_k_29);
	assign w_sys_tmp11743 = 32'sh00001691;
	assign w_sys_tmp11747 = (w_sys_tmp11748 + r_run_k_29);
	assign w_sys_tmp11748 = 32'sh000016f6;
	assign w_sys_tmp11752 = (w_sys_tmp11753 + r_run_k_29);
	assign w_sys_tmp11753 = 32'sh0000175b;
	assign w_sys_tmp11757 = (w_sys_tmp11758 + r_run_k_29);
	assign w_sys_tmp11758 = 32'sh000017c0;
	assign w_sys_tmp11762 = (w_sys_tmp11763 + r_run_k_29);
	assign w_sys_tmp11763 = 32'sh00001825;
	assign w_sys_tmp11767 = (w_sys_tmp11768 + r_run_k_29);
	assign w_sys_tmp11768 = 32'sh0000188a;
	assign w_sys_tmp11772 = (w_sys_tmp11773 + r_run_k_29);
	assign w_sys_tmp11773 = 32'sh000018ef;
	assign w_sys_tmp11777 = (w_sys_tmp11778 + r_run_k_29);
	assign w_sys_tmp11778 = 32'sh00001954;
	assign w_sys_tmp11782 = (w_sys_tmp11783 + r_run_k_29);
	assign w_sys_tmp11783 = 32'sh000019b9;
	assign w_sys_tmp11787 = (w_sys_tmp11788 + r_run_k_29);
	assign w_sys_tmp11788 = 32'sh00001a1e;
	assign w_sys_tmp11792 = (w_sys_tmp11793 + r_run_k_29);
	assign w_sys_tmp11793 = 32'sh00001a83;
	assign w_sys_tmp11797 = (w_sys_tmp11798 + r_run_k_29);
	assign w_sys_tmp11798 = 32'sh00001ae8;
	assign w_sys_tmp11802 = (w_sys_tmp11803 + r_run_k_29);
	assign w_sys_tmp11803 = 32'sh00001b4d;
	assign w_sys_tmp11807 = (w_sys_tmp11808 + r_run_k_29);
	assign w_sys_tmp11808 = 32'sh00001bb2;
	assign w_sys_tmp11812 = (w_sys_tmp11813 + r_run_k_29);
	assign w_sys_tmp11813 = 32'sh00001c17;
	assign w_sys_tmp11817 = (w_sys_tmp11818 + r_run_k_29);
	assign w_sys_tmp11818 = 32'sh00001c7c;
	assign w_sys_tmp11822 = (w_sys_tmp11823 + r_run_k_29);
	assign w_sys_tmp11823 = 32'sh00001ce1;
	assign w_sys_tmp11827 = (w_sys_tmp11828 + r_run_k_29);
	assign w_sys_tmp11828 = 32'sh00001d46;
	assign w_sys_tmp11832 = (w_sys_tmp11833 + r_run_k_29);
	assign w_sys_tmp11833 = 32'sh00001dab;
	assign w_sys_tmp11837 = (w_sys_tmp11838 + r_run_k_29);
	assign w_sys_tmp11838 = 32'sh00001e10;
	assign w_sys_tmp11842 = (w_sys_tmp11843 + r_run_k_29);
	assign w_sys_tmp11843 = 32'sh00001e75;
	assign w_sys_tmp11847 = (w_sys_tmp11848 + r_run_k_29);
	assign w_sys_tmp11848 = 32'sh00001eda;
	assign w_sys_tmp11852 = (w_sys_tmp11853 + r_run_k_29);
	assign w_sys_tmp11853 = 32'sh00001f3f;
	assign w_sys_tmp11857 = (w_sys_tmp11858 + r_run_k_29);
	assign w_sys_tmp11858 = 32'sh00001fa4;
	assign w_sys_tmp11862 = (w_sys_tmp11863 + r_run_k_29);
	assign w_sys_tmp11863 = 32'sh00002009;
	assign w_sys_tmp11867 = (w_sys_tmp11868 + r_run_k_29);
	assign w_sys_tmp11868 = 32'sh0000206e;
	assign w_sys_tmp11872 = (w_sys_tmp11873 + r_run_k_29);
	assign w_sys_tmp11873 = 32'sh000020d3;
	assign w_sys_tmp11877 = (w_sys_tmp11878 + r_run_k_29);
	assign w_sys_tmp11878 = 32'sh00002138;
	assign w_sys_tmp11882 = (w_sys_tmp11883 + r_run_k_29);
	assign w_sys_tmp11883 = 32'sh0000219d;
	assign w_sys_tmp11887 = (w_sys_tmp11888 + r_run_k_29);
	assign w_sys_tmp11888 = 32'sh00002202;
	assign w_sys_tmp11892 = (w_sys_tmp11893 + r_run_k_29);
	assign w_sys_tmp11893 = 32'sh00002267;
	assign w_sys_tmp11897 = (w_sys_tmp11898 + r_run_k_29);
	assign w_sys_tmp11898 = 32'sh000022cc;
	assign w_sys_tmp11902 = (w_sys_tmp11903 + r_run_k_29);
	assign w_sys_tmp11903 = 32'sh00002331;
	assign w_sys_tmp11907 = (w_sys_tmp11908 + r_run_k_29);
	assign w_sys_tmp11908 = 32'sh00002396;
	assign w_sys_tmp11912 = (w_sys_tmp11913 + r_run_k_29);
	assign w_sys_tmp11913 = 32'sh000023fb;
	assign w_sys_tmp11917 = (w_sys_tmp11918 + r_run_k_29);
	assign w_sys_tmp11918 = 32'sh00002460;
	assign w_sys_tmp11922 = (w_sys_tmp11923 + r_run_k_29);
	assign w_sys_tmp11923 = 32'sh000024c5;
	assign w_sys_tmp11927 = (w_sys_tmp11928 + r_run_k_29);
	assign w_sys_tmp11928 = 32'sh0000252a;
	assign w_sys_tmp11932 = (w_sys_tmp11933 + r_run_k_29);
	assign w_sys_tmp11933 = 32'sh0000258f;
	assign w_sys_tmp11937 = (w_sys_tmp11938 + r_run_k_29);
	assign w_sys_tmp11938 = 32'sh000025f4;
	assign w_sys_tmp11942 = (w_sys_tmp11943 + r_run_k_29);
	assign w_sys_tmp11943 = 32'sh00002659;
	assign w_sys_tmp11947 = (w_sys_tmp11948 + r_run_k_29);
	assign w_sys_tmp11948 = 32'sh000026be;
	assign w_sys_tmp11952 = (w_sys_tmp11953 + r_run_k_29);
	assign w_sys_tmp11953 = 32'sh00002723;
	assign w_sys_tmp11957 = (w_sys_tmp11958 + r_run_k_29);
	assign w_sys_tmp11958 = 32'sh00002788;
	assign w_sys_tmp11962 = (w_sys_tmp11963 + r_run_k_29);
	assign w_sys_tmp11963 = 32'sh000000f2;
	assign w_sys_tmp11967 = (w_sys_tmp11968 + r_run_k_29);
	assign w_sys_tmp11968 = 32'sh00000157;
	assign w_sys_tmp11972 = (w_sys_tmp11973 + r_run_k_29);
	assign w_sys_tmp11973 = 32'sh000001bc;
	assign w_sys_tmp11977 = (w_sys_tmp11978 + r_run_k_29);
	assign w_sys_tmp11978 = 32'sh00000221;
	assign w_sys_tmp11982 = (w_sys_tmp11983 + r_run_k_29);
	assign w_sys_tmp11983 = 32'sh00000286;
	assign w_sys_tmp11987 = (w_sys_tmp11988 + r_run_k_29);
	assign w_sys_tmp11988 = 32'sh000002eb;
	assign w_sys_tmp11992 = (w_sys_tmp11993 + r_run_k_29);
	assign w_sys_tmp11993 = 32'sh00000350;
	assign w_sys_tmp11997 = (w_sys_tmp11998 + r_run_k_29);
	assign w_sys_tmp11998 = 32'sh000003b5;
	assign w_sys_tmp12002 = (w_sys_tmp12003 + r_run_k_29);
	assign w_sys_tmp12003 = 32'sh0000041a;
	assign w_sys_tmp12007 = (w_sys_tmp12008 + r_run_k_29);
	assign w_sys_tmp12008 = 32'sh0000047f;
	assign w_sys_tmp12012 = (w_sys_tmp12013 + r_run_k_29);
	assign w_sys_tmp12013 = 32'sh000004e4;
	assign w_sys_tmp12017 = (w_sys_tmp12018 + r_run_k_29);
	assign w_sys_tmp12018 = 32'sh00000549;
	assign w_sys_tmp12022 = (w_sys_tmp12023 + r_run_k_29);
	assign w_sys_tmp12023 = 32'sh000005ae;
	assign w_sys_tmp12027 = (w_sys_tmp12028 + r_run_k_29);
	assign w_sys_tmp12028 = 32'sh00000613;
	assign w_sys_tmp12032 = (w_sys_tmp12033 + r_run_k_29);
	assign w_sys_tmp12033 = 32'sh00000678;
	assign w_sys_tmp12037 = (w_sys_tmp12038 + r_run_k_29);
	assign w_sys_tmp12038 = 32'sh000006dd;
	assign w_sys_tmp12042 = (w_sys_tmp12043 + r_run_k_29);
	assign w_sys_tmp12043 = 32'sh00000742;
	assign w_sys_tmp12047 = (w_sys_tmp12048 + r_run_k_29);
	assign w_sys_tmp12048 = 32'sh000007a7;
	assign w_sys_tmp12052 = (w_sys_tmp12053 + r_run_k_29);
	assign w_sys_tmp12053 = 32'sh0000080c;
	assign w_sys_tmp12057 = (w_sys_tmp12058 + r_run_k_29);
	assign w_sys_tmp12058 = 32'sh00000871;
	assign w_sys_tmp12062 = (w_sys_tmp12063 + r_run_k_29);
	assign w_sys_tmp12063 = 32'sh000008d6;
	assign w_sys_tmp12067 = (w_sys_tmp12068 + r_run_k_29);
	assign w_sys_tmp12068 = 32'sh0000093b;
	assign w_sys_tmp12072 = (w_sys_tmp12073 + r_run_k_29);
	assign w_sys_tmp12073 = 32'sh000009a0;
	assign w_sys_tmp12077 = (w_sys_tmp12078 + r_run_k_29);
	assign w_sys_tmp12078 = 32'sh00000a05;
	assign w_sys_tmp12082 = (w_sys_tmp12083 + r_run_k_29);
	assign w_sys_tmp12083 = 32'sh00000a6a;
	assign w_sys_tmp12087 = (w_sys_tmp12088 + r_run_k_29);
	assign w_sys_tmp12088 = 32'sh00000acf;
	assign w_sys_tmp12092 = (w_sys_tmp12093 + r_run_k_29);
	assign w_sys_tmp12093 = 32'sh00000b34;
	assign w_sys_tmp12097 = (w_sys_tmp12098 + r_run_k_29);
	assign w_sys_tmp12098 = 32'sh00000b99;
	assign w_sys_tmp12102 = (w_sys_tmp12103 + r_run_k_29);
	assign w_sys_tmp12103 = 32'sh00000bfe;
	assign w_sys_tmp12107 = (w_sys_tmp12108 + r_run_k_29);
	assign w_sys_tmp12108 = 32'sh00000c63;
	assign w_sys_tmp12112 = (w_sys_tmp12113 + r_run_k_29);
	assign w_sys_tmp12113 = 32'sh00000cc8;
	assign w_sys_tmp12117 = (w_sys_tmp12118 + r_run_k_29);
	assign w_sys_tmp12118 = 32'sh00000d2d;
	assign w_sys_tmp12122 = (w_sys_tmp12123 + r_run_k_29);
	assign w_sys_tmp12123 = 32'sh00000d92;
	assign w_sys_tmp12127 = (w_sys_tmp12128 + r_run_k_29);
	assign w_sys_tmp12128 = 32'sh00000df7;
	assign w_sys_tmp12132 = (w_sys_tmp12133 + r_run_k_29);
	assign w_sys_tmp12133 = 32'sh00000e5c;
	assign w_sys_tmp12137 = (w_sys_tmp12138 + r_run_k_29);
	assign w_sys_tmp12138 = 32'sh00000ec1;
	assign w_sys_tmp12142 = (w_sys_tmp12143 + r_run_k_29);
	assign w_sys_tmp12143 = 32'sh00000f26;
	assign w_sys_tmp12147 = (w_sys_tmp12148 + r_run_k_29);
	assign w_sys_tmp12148 = 32'sh00000f8b;
	assign w_sys_tmp12152 = (w_sys_tmp12153 + r_run_k_29);
	assign w_sys_tmp12153 = 32'sh00000ff0;
	assign w_sys_tmp12157 = (w_sys_tmp12158 + r_run_k_29);
	assign w_sys_tmp12158 = 32'sh00001055;
	assign w_sys_tmp12162 = (w_sys_tmp12163 + r_run_k_29);
	assign w_sys_tmp12163 = 32'sh000010ba;
	assign w_sys_tmp12167 = (w_sys_tmp12168 + r_run_k_29);
	assign w_sys_tmp12168 = 32'sh0000111f;
	assign w_sys_tmp12172 = (w_sys_tmp12173 + r_run_k_29);
	assign w_sys_tmp12173 = 32'sh00001184;
	assign w_sys_tmp12177 = (w_sys_tmp12178 + r_run_k_29);
	assign w_sys_tmp12178 = 32'sh000011e9;
	assign w_sys_tmp12182 = (w_sys_tmp12183 + r_run_k_29);
	assign w_sys_tmp12183 = 32'sh0000124e;
	assign w_sys_tmp12187 = (w_sys_tmp12188 + r_run_k_29);
	assign w_sys_tmp12188 = 32'sh000012b3;
	assign w_sys_tmp12192 = (w_sys_tmp12193 + r_run_k_29);
	assign w_sys_tmp12193 = 32'sh00001318;
	assign w_sys_tmp12197 = (w_sys_tmp12198 + r_run_k_29);
	assign w_sys_tmp12198 = 32'sh0000137d;
	assign w_sys_tmp12202 = (w_sys_tmp12203 + r_run_k_29);
	assign w_sys_tmp12203 = 32'sh000013e2;
	assign w_sys_tmp12207 = (w_sys_tmp12208 + r_run_k_29);
	assign w_sys_tmp12208 = 32'sh00001447;
	assign w_sys_tmp12212 = (w_sys_tmp12213 + r_run_k_29);
	assign w_sys_tmp12213 = 32'sh000014ac;
	assign w_sys_tmp12217 = (w_sys_tmp12218 + r_run_k_29);
	assign w_sys_tmp12218 = 32'sh00001511;
	assign w_sys_tmp12222 = (w_sys_tmp12223 + r_run_k_29);
	assign w_sys_tmp12223 = 32'sh00001576;
	assign w_sys_tmp12227 = (w_sys_tmp12228 + r_run_k_29);
	assign w_sys_tmp12228 = 32'sh000015db;
	assign w_sys_tmp12232 = (w_sys_tmp12233 + r_run_k_29);
	assign w_sys_tmp12233 = 32'sh00001640;
	assign w_sys_tmp12237 = (w_sys_tmp12238 + r_run_k_29);
	assign w_sys_tmp12238 = 32'sh000016a5;
	assign w_sys_tmp12242 = (w_sys_tmp12243 + r_run_k_29);
	assign w_sys_tmp12243 = 32'sh0000170a;
	assign w_sys_tmp12247 = (w_sys_tmp12248 + r_run_k_29);
	assign w_sys_tmp12248 = 32'sh0000176f;
	assign w_sys_tmp12252 = (w_sys_tmp12253 + r_run_k_29);
	assign w_sys_tmp12253 = 32'sh000017d4;
	assign w_sys_tmp12257 = (w_sys_tmp12258 + r_run_k_29);
	assign w_sys_tmp12258 = 32'sh00001839;
	assign w_sys_tmp12262 = (w_sys_tmp12263 + r_run_k_29);
	assign w_sys_tmp12263 = 32'sh0000189e;
	assign w_sys_tmp12267 = (w_sys_tmp12268 + r_run_k_29);
	assign w_sys_tmp12268 = 32'sh00001903;
	assign w_sys_tmp12272 = (w_sys_tmp12273 + r_run_k_29);
	assign w_sys_tmp12273 = 32'sh00001968;
	assign w_sys_tmp12277 = (w_sys_tmp12278 + r_run_k_29);
	assign w_sys_tmp12278 = 32'sh000019cd;
	assign w_sys_tmp12282 = (w_sys_tmp12283 + r_run_k_29);
	assign w_sys_tmp12283 = 32'sh00001a32;
	assign w_sys_tmp12287 = (w_sys_tmp12288 + r_run_k_29);
	assign w_sys_tmp12288 = 32'sh00001a97;
	assign w_sys_tmp12292 = (w_sys_tmp12293 + r_run_k_29);
	assign w_sys_tmp12293 = 32'sh00001afc;
	assign w_sys_tmp12297 = (w_sys_tmp12298 + r_run_k_29);
	assign w_sys_tmp12298 = 32'sh00001b61;
	assign w_sys_tmp12302 = (w_sys_tmp12303 + r_run_k_29);
	assign w_sys_tmp12303 = 32'sh00001bc6;
	assign w_sys_tmp12307 = (w_sys_tmp12308 + r_run_k_29);
	assign w_sys_tmp12308 = 32'sh00001c2b;
	assign w_sys_tmp12312 = (w_sys_tmp12313 + r_run_k_29);
	assign w_sys_tmp12313 = 32'sh00001c90;
	assign w_sys_tmp12317 = (w_sys_tmp12318 + r_run_k_29);
	assign w_sys_tmp12318 = 32'sh00001cf5;
	assign w_sys_tmp12322 = (w_sys_tmp12323 + r_run_k_29);
	assign w_sys_tmp12323 = 32'sh00001d5a;
	assign w_sys_tmp12327 = (w_sys_tmp12328 + r_run_k_29);
	assign w_sys_tmp12328 = 32'sh00001dbf;
	assign w_sys_tmp12332 = (w_sys_tmp12333 + r_run_k_29);
	assign w_sys_tmp12333 = 32'sh00001e24;
	assign w_sys_tmp12337 = (w_sys_tmp12338 + r_run_k_29);
	assign w_sys_tmp12338 = 32'sh00001e89;
	assign w_sys_tmp12342 = (w_sys_tmp12343 + r_run_k_29);
	assign w_sys_tmp12343 = 32'sh00001eee;
	assign w_sys_tmp12347 = (w_sys_tmp12348 + r_run_k_29);
	assign w_sys_tmp12348 = 32'sh00001f53;
	assign w_sys_tmp12352 = (w_sys_tmp12353 + r_run_k_29);
	assign w_sys_tmp12353 = 32'sh00001fb8;
	assign w_sys_tmp12357 = (w_sys_tmp12358 + r_run_k_29);
	assign w_sys_tmp12358 = 32'sh0000201d;
	assign w_sys_tmp12362 = (w_sys_tmp12363 + r_run_k_29);
	assign w_sys_tmp12363 = 32'sh00002082;
	assign w_sys_tmp12367 = (w_sys_tmp12368 + r_run_k_29);
	assign w_sys_tmp12368 = 32'sh000020e7;
	assign w_sys_tmp12372 = (w_sys_tmp12373 + r_run_k_29);
	assign w_sys_tmp12373 = 32'sh0000214c;
	assign w_sys_tmp12377 = (w_sys_tmp12378 + r_run_k_29);
	assign w_sys_tmp12378 = 32'sh000021b1;
	assign w_sys_tmp12382 = (w_sys_tmp12383 + r_run_k_29);
	assign w_sys_tmp12383 = 32'sh00002216;
	assign w_sys_tmp12387 = (w_sys_tmp12388 + r_run_k_29);
	assign w_sys_tmp12388 = 32'sh0000227b;
	assign w_sys_tmp12392 = (w_sys_tmp12393 + r_run_k_29);
	assign w_sys_tmp12393 = 32'sh000022e0;
	assign w_sys_tmp12397 = (w_sys_tmp12398 + r_run_k_29);
	assign w_sys_tmp12398 = 32'sh00002345;
	assign w_sys_tmp12402 = (w_sys_tmp12403 + r_run_k_29);
	assign w_sys_tmp12403 = 32'sh000023aa;
	assign w_sys_tmp12407 = (w_sys_tmp12408 + r_run_k_29);
	assign w_sys_tmp12408 = 32'sh0000240f;
	assign w_sys_tmp12412 = (w_sys_tmp12413 + r_run_k_29);
	assign w_sys_tmp12413 = 32'sh00002474;
	assign w_sys_tmp12417 = (w_sys_tmp12418 + r_run_k_29);
	assign w_sys_tmp12418 = 32'sh000024d9;
	assign w_sys_tmp12422 = (w_sys_tmp12423 + r_run_k_29);
	assign w_sys_tmp12423 = 32'sh0000253e;
	assign w_sys_tmp12427 = (w_sys_tmp12428 + r_run_k_29);
	assign w_sys_tmp12428 = 32'sh000025a3;
	assign w_sys_tmp12432 = (w_sys_tmp12433 + r_run_k_29);
	assign w_sys_tmp12433 = 32'sh00002608;
	assign w_sys_tmp12437 = (w_sys_tmp12438 + r_run_k_29);
	assign w_sys_tmp12438 = 32'sh0000266d;
	assign w_sys_tmp12442 = (w_sys_tmp12443 + r_run_k_29);
	assign w_sys_tmp12443 = 32'sh000026d2;
	assign w_sys_tmp12447 = (w_sys_tmp12448 + r_run_k_29);
	assign w_sys_tmp12448 = 32'sh00002737;
	assign w_sys_tmp12452 = (w_sys_tmp12453 + r_run_k_29);
	assign w_sys_tmp12453 = 32'sh0000279c;
	assign w_sys_tmp12457 = (w_sys_tmp12458 + r_run_k_29);
	assign w_sys_tmp12458 = 32'sh00000106;
	assign w_sys_tmp12462 = (w_sys_tmp12463 + r_run_k_29);
	assign w_sys_tmp12463 = 32'sh0000016b;
	assign w_sys_tmp12467 = (w_sys_tmp12468 + r_run_k_29);
	assign w_sys_tmp12468 = 32'sh000001d0;
	assign w_sys_tmp12472 = (w_sys_tmp12473 + r_run_k_29);
	assign w_sys_tmp12473 = 32'sh00000235;
	assign w_sys_tmp12477 = (w_sys_tmp12478 + r_run_k_29);
	assign w_sys_tmp12478 = 32'sh0000029a;
	assign w_sys_tmp12482 = (w_sys_tmp12483 + r_run_k_29);
	assign w_sys_tmp12483 = 32'sh000002ff;
	assign w_sys_tmp12487 = (w_sys_tmp12488 + r_run_k_29);
	assign w_sys_tmp12488 = 32'sh00000364;
	assign w_sys_tmp12492 = (w_sys_tmp12493 + r_run_k_29);
	assign w_sys_tmp12493 = 32'sh000003c9;
	assign w_sys_tmp12497 = (w_sys_tmp12498 + r_run_k_29);
	assign w_sys_tmp12498 = 32'sh0000042e;
	assign w_sys_tmp12502 = (w_sys_tmp12503 + r_run_k_29);
	assign w_sys_tmp12503 = 32'sh00000493;
	assign w_sys_tmp12507 = (w_sys_tmp12508 + r_run_k_29);
	assign w_sys_tmp12508 = 32'sh000004f8;
	assign w_sys_tmp12512 = (w_sys_tmp12513 + r_run_k_29);
	assign w_sys_tmp12513 = 32'sh0000055d;
	assign w_sys_tmp12517 = (w_sys_tmp12518 + r_run_k_29);
	assign w_sys_tmp12518 = 32'sh000005c2;
	assign w_sys_tmp12522 = (w_sys_tmp12523 + r_run_k_29);
	assign w_sys_tmp12523 = 32'sh00000627;
	assign w_sys_tmp12527 = (w_sys_tmp12528 + r_run_k_29);
	assign w_sys_tmp12528 = 32'sh0000068c;
	assign w_sys_tmp12532 = (w_sys_tmp12533 + r_run_k_29);
	assign w_sys_tmp12533 = 32'sh000006f1;
	assign w_sys_tmp12537 = (w_sys_tmp12538 + r_run_k_29);
	assign w_sys_tmp12538 = 32'sh00000756;
	assign w_sys_tmp12542 = (w_sys_tmp12543 + r_run_k_29);
	assign w_sys_tmp12543 = 32'sh000007bb;
	assign w_sys_tmp12547 = (w_sys_tmp12548 + r_run_k_29);
	assign w_sys_tmp12548 = 32'sh00000820;
	assign w_sys_tmp12552 = (w_sys_tmp12553 + r_run_k_29);
	assign w_sys_tmp12553 = 32'sh00000885;
	assign w_sys_tmp12557 = (w_sys_tmp12558 + r_run_k_29);
	assign w_sys_tmp12558 = 32'sh000008ea;
	assign w_sys_tmp12562 = (w_sys_tmp12563 + r_run_k_29);
	assign w_sys_tmp12563 = 32'sh0000094f;
	assign w_sys_tmp12567 = (w_sys_tmp12568 + r_run_k_29);
	assign w_sys_tmp12568 = 32'sh000009b4;
	assign w_sys_tmp12572 = (w_sys_tmp12573 + r_run_k_29);
	assign w_sys_tmp12573 = 32'sh00000a19;
	assign w_sys_tmp12577 = (w_sys_tmp12578 + r_run_k_29);
	assign w_sys_tmp12578 = 32'sh00000a7e;
	assign w_sys_tmp12582 = (w_sys_tmp12583 + r_run_k_29);
	assign w_sys_tmp12583 = 32'sh00000ae3;
	assign w_sys_tmp12587 = (w_sys_tmp12588 + r_run_k_29);
	assign w_sys_tmp12588 = 32'sh00000b48;
	assign w_sys_tmp12592 = (w_sys_tmp12593 + r_run_k_29);
	assign w_sys_tmp12593 = 32'sh00000bad;
	assign w_sys_tmp12597 = (w_sys_tmp12598 + r_run_k_29);
	assign w_sys_tmp12598 = 32'sh00000c12;
	assign w_sys_tmp12602 = (w_sys_tmp12603 + r_run_k_29);
	assign w_sys_tmp12603 = 32'sh00000c77;
	assign w_sys_tmp12607 = (w_sys_tmp12608 + r_run_k_29);
	assign w_sys_tmp12608 = 32'sh00000cdc;
	assign w_sys_tmp12612 = (w_sys_tmp12613 + r_run_k_29);
	assign w_sys_tmp12613 = 32'sh00000d41;
	assign w_sys_tmp12617 = (w_sys_tmp12618 + r_run_k_29);
	assign w_sys_tmp12618 = 32'sh00000da6;
	assign w_sys_tmp12622 = (w_sys_tmp12623 + r_run_k_29);
	assign w_sys_tmp12623 = 32'sh00000e0b;
	assign w_sys_tmp12627 = (w_sys_tmp12628 + r_run_k_29);
	assign w_sys_tmp12628 = 32'sh00000e70;
	assign w_sys_tmp12632 = (w_sys_tmp12633 + r_run_k_29);
	assign w_sys_tmp12633 = 32'sh00000ed5;
	assign w_sys_tmp12637 = (w_sys_tmp12638 + r_run_k_29);
	assign w_sys_tmp12638 = 32'sh00000f3a;
	assign w_sys_tmp12642 = (w_sys_tmp12643 + r_run_k_29);
	assign w_sys_tmp12643 = 32'sh00000f9f;
	assign w_sys_tmp12647 = (w_sys_tmp12648 + r_run_k_29);
	assign w_sys_tmp12648 = 32'sh00001004;
	assign w_sys_tmp12652 = (w_sys_tmp12653 + r_run_k_29);
	assign w_sys_tmp12653 = 32'sh00001069;
	assign w_sys_tmp12657 = (w_sys_tmp12658 + r_run_k_29);
	assign w_sys_tmp12658 = 32'sh000010ce;
	assign w_sys_tmp12662 = (w_sys_tmp12663 + r_run_k_29);
	assign w_sys_tmp12663 = 32'sh00001133;
	assign w_sys_tmp12667 = (w_sys_tmp12668 + r_run_k_29);
	assign w_sys_tmp12668 = 32'sh00001198;
	assign w_sys_tmp12672 = (w_sys_tmp12673 + r_run_k_29);
	assign w_sys_tmp12673 = 32'sh000011fd;
	assign w_sys_tmp12677 = (w_sys_tmp12678 + r_run_k_29);
	assign w_sys_tmp12678 = 32'sh00001262;
	assign w_sys_tmp12682 = (w_sys_tmp12683 + r_run_k_29);
	assign w_sys_tmp12683 = 32'sh000012c7;
	assign w_sys_tmp12687 = (w_sys_tmp12688 + r_run_k_29);
	assign w_sys_tmp12688 = 32'sh0000132c;
	assign w_sys_tmp12692 = (w_sys_tmp12693 + r_run_k_29);
	assign w_sys_tmp12693 = 32'sh00001391;
	assign w_sys_tmp12697 = (w_sys_tmp12698 + r_run_k_29);
	assign w_sys_tmp12698 = 32'sh000013f6;
	assign w_sys_tmp12702 = (w_sys_tmp12703 + r_run_k_29);
	assign w_sys_tmp12703 = 32'sh0000145b;
	assign w_sys_tmp12707 = (w_sys_tmp12708 + r_run_k_29);
	assign w_sys_tmp12708 = 32'sh000014c0;
	assign w_sys_tmp12712 = (w_sys_tmp12713 + r_run_k_29);
	assign w_sys_tmp12713 = 32'sh00001525;
	assign w_sys_tmp12717 = (w_sys_tmp12718 + r_run_k_29);
	assign w_sys_tmp12718 = 32'sh0000158a;
	assign w_sys_tmp12722 = (w_sys_tmp12723 + r_run_k_29);
	assign w_sys_tmp12723 = 32'sh000015ef;
	assign w_sys_tmp12727 = (w_sys_tmp12728 + r_run_k_29);
	assign w_sys_tmp12728 = 32'sh00001654;
	assign w_sys_tmp12732 = (w_sys_tmp12733 + r_run_k_29);
	assign w_sys_tmp12733 = 32'sh000016b9;
	assign w_sys_tmp12737 = (w_sys_tmp12738 + r_run_k_29);
	assign w_sys_tmp12738 = 32'sh0000171e;
	assign w_sys_tmp12742 = (w_sys_tmp12743 + r_run_k_29);
	assign w_sys_tmp12743 = 32'sh00001783;
	assign w_sys_tmp12747 = (w_sys_tmp12748 + r_run_k_29);
	assign w_sys_tmp12748 = 32'sh000017e8;
	assign w_sys_tmp12752 = (w_sys_tmp12753 + r_run_k_29);
	assign w_sys_tmp12753 = 32'sh0000184d;
	assign w_sys_tmp12757 = (w_sys_tmp12758 + r_run_k_29);
	assign w_sys_tmp12758 = 32'sh000018b2;
	assign w_sys_tmp12762 = (w_sys_tmp12763 + r_run_k_29);
	assign w_sys_tmp12763 = 32'sh00001917;
	assign w_sys_tmp12767 = (w_sys_tmp12768 + r_run_k_29);
	assign w_sys_tmp12768 = 32'sh0000197c;
	assign w_sys_tmp12772 = (w_sys_tmp12773 + r_run_k_29);
	assign w_sys_tmp12773 = 32'sh000019e1;
	assign w_sys_tmp12777 = (w_sys_tmp12778 + r_run_k_29);
	assign w_sys_tmp12778 = 32'sh00001a46;
	assign w_sys_tmp12782 = (w_sys_tmp12783 + r_run_k_29);
	assign w_sys_tmp12783 = 32'sh00001aab;
	assign w_sys_tmp12787 = (w_sys_tmp12788 + r_run_k_29);
	assign w_sys_tmp12788 = 32'sh00001b10;
	assign w_sys_tmp12792 = (w_sys_tmp12793 + r_run_k_29);
	assign w_sys_tmp12793 = 32'sh00001b75;
	assign w_sys_tmp12797 = (w_sys_tmp12798 + r_run_k_29);
	assign w_sys_tmp12798 = 32'sh00001bda;
	assign w_sys_tmp12802 = (w_sys_tmp12803 + r_run_k_29);
	assign w_sys_tmp12803 = 32'sh00001c3f;
	assign w_sys_tmp12807 = (w_sys_tmp12808 + r_run_k_29);
	assign w_sys_tmp12808 = 32'sh00001ca4;
	assign w_sys_tmp12812 = (w_sys_tmp12813 + r_run_k_29);
	assign w_sys_tmp12813 = 32'sh00001d09;
	assign w_sys_tmp12817 = (w_sys_tmp12818 + r_run_k_29);
	assign w_sys_tmp12818 = 32'sh00001d6e;
	assign w_sys_tmp12822 = (w_sys_tmp12823 + r_run_k_29);
	assign w_sys_tmp12823 = 32'sh00001dd3;
	assign w_sys_tmp12827 = (w_sys_tmp12828 + r_run_k_29);
	assign w_sys_tmp12828 = 32'sh00001e38;
	assign w_sys_tmp12832 = (w_sys_tmp12833 + r_run_k_29);
	assign w_sys_tmp12833 = 32'sh00001e9d;
	assign w_sys_tmp12837 = (w_sys_tmp12838 + r_run_k_29);
	assign w_sys_tmp12838 = 32'sh00001f02;
	assign w_sys_tmp12842 = (w_sys_tmp12843 + r_run_k_29);
	assign w_sys_tmp12843 = 32'sh00001f67;
	assign w_sys_tmp12847 = (w_sys_tmp12848 + r_run_k_29);
	assign w_sys_tmp12848 = 32'sh00001fcc;
	assign w_sys_tmp12852 = (w_sys_tmp12853 + r_run_k_29);
	assign w_sys_tmp12853 = 32'sh00002031;
	assign w_sys_tmp12857 = (w_sys_tmp12858 + r_run_k_29);
	assign w_sys_tmp12858 = 32'sh00002096;
	assign w_sys_tmp12862 = (w_sys_tmp12863 + r_run_k_29);
	assign w_sys_tmp12863 = 32'sh000020fb;
	assign w_sys_tmp12867 = (w_sys_tmp12868 + r_run_k_29);
	assign w_sys_tmp12868 = 32'sh00002160;
	assign w_sys_tmp12872 = (w_sys_tmp12873 + r_run_k_29);
	assign w_sys_tmp12873 = 32'sh000021c5;
	assign w_sys_tmp12877 = (w_sys_tmp12878 + r_run_k_29);
	assign w_sys_tmp12878 = 32'sh0000222a;
	assign w_sys_tmp12882 = (w_sys_tmp12883 + r_run_k_29);
	assign w_sys_tmp12883 = 32'sh0000228f;
	assign w_sys_tmp12887 = (w_sys_tmp12888 + r_run_k_29);
	assign w_sys_tmp12888 = 32'sh000022f4;
	assign w_sys_tmp12892 = (w_sys_tmp12893 + r_run_k_29);
	assign w_sys_tmp12893 = 32'sh00002359;
	assign w_sys_tmp12897 = (w_sys_tmp12898 + r_run_k_29);
	assign w_sys_tmp12898 = 32'sh000023be;
	assign w_sys_tmp12902 = (w_sys_tmp12903 + r_run_k_29);
	assign w_sys_tmp12903 = 32'sh00002423;
	assign w_sys_tmp12907 = (w_sys_tmp12908 + r_run_k_29);
	assign w_sys_tmp12908 = 32'sh00002488;
	assign w_sys_tmp12912 = (w_sys_tmp12913 + r_run_k_29);
	assign w_sys_tmp12913 = 32'sh000024ed;
	assign w_sys_tmp12917 = (w_sys_tmp12918 + r_run_k_29);
	assign w_sys_tmp12918 = 32'sh00002552;
	assign w_sys_tmp12922 = (w_sys_tmp12923 + r_run_k_29);
	assign w_sys_tmp12923 = 32'sh000025b7;
	assign w_sys_tmp12927 = (w_sys_tmp12928 + r_run_k_29);
	assign w_sys_tmp12928 = 32'sh0000261c;
	assign w_sys_tmp12932 = (w_sys_tmp12933 + r_run_k_29);
	assign w_sys_tmp12933 = 32'sh00002681;
	assign w_sys_tmp12937 = (w_sys_tmp12938 + r_run_k_29);
	assign w_sys_tmp12938 = 32'sh000026e6;
	assign w_sys_tmp12942 = (w_sys_tmp12943 + r_run_k_29);
	assign w_sys_tmp12943 = 32'sh0000274b;
	assign w_sys_tmp12947 = (w_sys_tmp12948 + r_run_k_29);
	assign w_sys_tmp12948 = 32'sh000027b0;
	assign w_sys_tmp12951 = (r_run_k_29 + w_sys_intOne);
	assign w_sys_tmp12952 = 32'sh0000001a;
	assign w_sys_tmp12953 = ( !w_sys_tmp12954 );
	assign w_sys_tmp12954 = (w_sys_tmp12955 < r_run_k_29);
	assign w_sys_tmp12955 = 32'sh0000001e;
	assign w_sys_tmp12958 = (w_sys_tmp12959 + r_run_k_29);
	assign w_sys_tmp12959 = 32'sh000000ca;
	assign w_sys_tmp12960 = w_sub20_result_dataout;
	assign w_sys_tmp12964 = (w_sys_tmp12965 + r_run_k_29);
	assign w_sys_tmp12965 = 32'sh0000012f;
	assign w_sys_tmp12970 = (w_sys_tmp12971 + r_run_k_29);
	assign w_sys_tmp12971 = 32'sh00000194;
	assign w_sys_tmp12976 = (w_sys_tmp12977 + r_run_k_29);
	assign w_sys_tmp12977 = 32'sh000001f9;
	assign w_sys_tmp12982 = (w_sys_tmp12983 + r_run_k_29);
	assign w_sys_tmp12983 = 32'sh0000025e;
	assign w_sys_tmp12988 = (w_sys_tmp12989 + r_run_k_29);
	assign w_sys_tmp12989 = 32'sh000002c3;
	assign w_sys_tmp12994 = (w_sys_tmp12995 + r_run_k_29);
	assign w_sys_tmp12995 = 32'sh00000328;
	assign w_sys_tmp13000 = (w_sys_tmp13001 + r_run_k_29);
	assign w_sys_tmp13001 = 32'sh0000038d;
	assign w_sys_tmp13006 = (w_sys_tmp13007 + r_run_k_29);
	assign w_sys_tmp13007 = 32'sh000003f2;
	assign w_sys_tmp13012 = (w_sys_tmp13013 + r_run_k_29);
	assign w_sys_tmp13013 = 32'sh00000457;
	assign w_sys_tmp13018 = (w_sys_tmp13019 + r_run_k_29);
	assign w_sys_tmp13019 = 32'sh000004bc;
	assign w_sys_tmp13024 = (w_sys_tmp13025 + r_run_k_29);
	assign w_sys_tmp13025 = 32'sh00000521;
	assign w_sys_tmp13030 = (w_sys_tmp13031 + r_run_k_29);
	assign w_sys_tmp13031 = 32'sh00000586;
	assign w_sys_tmp13036 = (w_sys_tmp13037 + r_run_k_29);
	assign w_sys_tmp13037 = 32'sh000005eb;
	assign w_sys_tmp13042 = (w_sys_tmp13043 + r_run_k_29);
	assign w_sys_tmp13043 = 32'sh00000650;
	assign w_sys_tmp13048 = (w_sys_tmp13049 + r_run_k_29);
	assign w_sys_tmp13049 = 32'sh000006b5;
	assign w_sys_tmp13054 = (w_sys_tmp13055 + r_run_k_29);
	assign w_sys_tmp13055 = 32'sh0000071a;
	assign w_sys_tmp13060 = (w_sys_tmp13061 + r_run_k_29);
	assign w_sys_tmp13061 = 32'sh0000077f;
	assign w_sys_tmp13066 = (w_sys_tmp13067 + r_run_k_29);
	assign w_sys_tmp13067 = 32'sh000007e4;
	assign w_sys_tmp13072 = (w_sys_tmp13073 + r_run_k_29);
	assign w_sys_tmp13073 = 32'sh00000849;
	assign w_sys_tmp13078 = (w_sys_tmp13079 + r_run_k_29);
	assign w_sys_tmp13079 = 32'sh000008ae;
	assign w_sys_tmp13083 = (w_sys_tmp13084 + r_run_k_29);
	assign w_sys_tmp13084 = 32'sh00000913;
	assign w_sys_tmp13088 = (w_sys_tmp13089 + r_run_k_29);
	assign w_sys_tmp13089 = 32'sh00000978;
	assign w_sys_tmp13093 = (w_sys_tmp13094 + r_run_k_29);
	assign w_sys_tmp13094 = 32'sh000009dd;
	assign w_sys_tmp13098 = (w_sys_tmp13099 + r_run_k_29);
	assign w_sys_tmp13099 = 32'sh00000a42;
	assign w_sys_tmp13103 = (w_sys_tmp13104 + r_run_k_29);
	assign w_sys_tmp13104 = 32'sh00000aa7;
	assign w_sys_tmp13108 = (w_sys_tmp13109 + r_run_k_29);
	assign w_sys_tmp13109 = 32'sh00000b0c;
	assign w_sys_tmp13113 = (w_sys_tmp13114 + r_run_k_29);
	assign w_sys_tmp13114 = 32'sh00000b71;
	assign w_sys_tmp13118 = (w_sys_tmp13119 + r_run_k_29);
	assign w_sys_tmp13119 = 32'sh00000bd6;
	assign w_sys_tmp13123 = (w_sys_tmp13124 + r_run_k_29);
	assign w_sys_tmp13124 = 32'sh00000c3b;
	assign w_sys_tmp13128 = (w_sys_tmp13129 + r_run_k_29);
	assign w_sys_tmp13129 = 32'sh00000ca0;
	assign w_sys_tmp13133 = (w_sys_tmp13134 + r_run_k_29);
	assign w_sys_tmp13134 = 32'sh00000d05;
	assign w_sys_tmp13138 = (w_sys_tmp13139 + r_run_k_29);
	assign w_sys_tmp13139 = 32'sh00000d6a;
	assign w_sys_tmp13143 = (w_sys_tmp13144 + r_run_k_29);
	assign w_sys_tmp13144 = 32'sh00000dcf;
	assign w_sys_tmp13148 = (w_sys_tmp13149 + r_run_k_29);
	assign w_sys_tmp13149 = 32'sh00000e34;
	assign w_sys_tmp13153 = (w_sys_tmp13154 + r_run_k_29);
	assign w_sys_tmp13154 = 32'sh00000e99;
	assign w_sys_tmp13158 = (w_sys_tmp13159 + r_run_k_29);
	assign w_sys_tmp13159 = 32'sh00000efe;
	assign w_sys_tmp13163 = (w_sys_tmp13164 + r_run_k_29);
	assign w_sys_tmp13164 = 32'sh00000f63;
	assign w_sys_tmp13168 = (w_sys_tmp13169 + r_run_k_29);
	assign w_sys_tmp13169 = 32'sh00000fc8;
	assign w_sys_tmp13173 = (w_sys_tmp13174 + r_run_k_29);
	assign w_sys_tmp13174 = 32'sh0000102d;
	assign w_sys_tmp13178 = (w_sys_tmp13179 + r_run_k_29);
	assign w_sys_tmp13179 = 32'sh00001092;
	assign w_sys_tmp13183 = (w_sys_tmp13184 + r_run_k_29);
	assign w_sys_tmp13184 = 32'sh000010f7;
	assign w_sys_tmp13188 = (w_sys_tmp13189 + r_run_k_29);
	assign w_sys_tmp13189 = 32'sh0000115c;
	assign w_sys_tmp13193 = (w_sys_tmp13194 + r_run_k_29);
	assign w_sys_tmp13194 = 32'sh000011c1;
	assign w_sys_tmp13198 = (w_sys_tmp13199 + r_run_k_29);
	assign w_sys_tmp13199 = 32'sh00001226;
	assign w_sys_tmp13203 = (w_sys_tmp13204 + r_run_k_29);
	assign w_sys_tmp13204 = 32'sh0000128b;
	assign w_sys_tmp13208 = (w_sys_tmp13209 + r_run_k_29);
	assign w_sys_tmp13209 = 32'sh000012f0;
	assign w_sys_tmp13213 = (w_sys_tmp13214 + r_run_k_29);
	assign w_sys_tmp13214 = 32'sh00001355;
	assign w_sys_tmp13218 = (w_sys_tmp13219 + r_run_k_29);
	assign w_sys_tmp13219 = 32'sh000013ba;
	assign w_sys_tmp13223 = (w_sys_tmp13224 + r_run_k_29);
	assign w_sys_tmp13224 = 32'sh0000141f;
	assign w_sys_tmp13228 = (w_sys_tmp13229 + r_run_k_29);
	assign w_sys_tmp13229 = 32'sh00001484;
	assign w_sys_tmp13233 = (w_sys_tmp13234 + r_run_k_29);
	assign w_sys_tmp13234 = 32'sh000014e9;
	assign w_sys_tmp13238 = (w_sys_tmp13239 + r_run_k_29);
	assign w_sys_tmp13239 = 32'sh0000154e;
	assign w_sys_tmp13243 = (w_sys_tmp13244 + r_run_k_29);
	assign w_sys_tmp13244 = 32'sh000015b3;
	assign w_sys_tmp13248 = (w_sys_tmp13249 + r_run_k_29);
	assign w_sys_tmp13249 = 32'sh00001618;
	assign w_sys_tmp13253 = (w_sys_tmp13254 + r_run_k_29);
	assign w_sys_tmp13254 = 32'sh0000167d;
	assign w_sys_tmp13258 = (w_sys_tmp13259 + r_run_k_29);
	assign w_sys_tmp13259 = 32'sh000016e2;
	assign w_sys_tmp13263 = (w_sys_tmp13264 + r_run_k_29);
	assign w_sys_tmp13264 = 32'sh00001747;
	assign w_sys_tmp13268 = (w_sys_tmp13269 + r_run_k_29);
	assign w_sys_tmp13269 = 32'sh000017ac;
	assign w_sys_tmp13273 = (w_sys_tmp13274 + r_run_k_29);
	assign w_sys_tmp13274 = 32'sh00001811;
	assign w_sys_tmp13278 = (w_sys_tmp13279 + r_run_k_29);
	assign w_sys_tmp13279 = 32'sh00001876;
	assign w_sys_tmp13283 = (w_sys_tmp13284 + r_run_k_29);
	assign w_sys_tmp13284 = 32'sh000018db;
	assign w_sys_tmp13288 = (w_sys_tmp13289 + r_run_k_29);
	assign w_sys_tmp13289 = 32'sh00001940;
	assign w_sys_tmp13293 = (w_sys_tmp13294 + r_run_k_29);
	assign w_sys_tmp13294 = 32'sh000019a5;
	assign w_sys_tmp13298 = (w_sys_tmp13299 + r_run_k_29);
	assign w_sys_tmp13299 = 32'sh00001a0a;
	assign w_sys_tmp13303 = (w_sys_tmp13304 + r_run_k_29);
	assign w_sys_tmp13304 = 32'sh00001a6f;
	assign w_sys_tmp13308 = (w_sys_tmp13309 + r_run_k_29);
	assign w_sys_tmp13309 = 32'sh00001ad4;
	assign w_sys_tmp13313 = (w_sys_tmp13314 + r_run_k_29);
	assign w_sys_tmp13314 = 32'sh00001b39;
	assign w_sys_tmp13318 = (w_sys_tmp13319 + r_run_k_29);
	assign w_sys_tmp13319 = 32'sh00001b9e;
	assign w_sys_tmp13323 = (w_sys_tmp13324 + r_run_k_29);
	assign w_sys_tmp13324 = 32'sh00001c03;
	assign w_sys_tmp13328 = (w_sys_tmp13329 + r_run_k_29);
	assign w_sys_tmp13329 = 32'sh00001c68;
	assign w_sys_tmp13333 = (w_sys_tmp13334 + r_run_k_29);
	assign w_sys_tmp13334 = 32'sh00001ccd;
	assign w_sys_tmp13338 = (w_sys_tmp13339 + r_run_k_29);
	assign w_sys_tmp13339 = 32'sh00001d32;
	assign w_sys_tmp13343 = (w_sys_tmp13344 + r_run_k_29);
	assign w_sys_tmp13344 = 32'sh00001d97;
	assign w_sys_tmp13348 = (w_sys_tmp13349 + r_run_k_29);
	assign w_sys_tmp13349 = 32'sh00001dfc;
	assign w_sys_tmp13353 = (w_sys_tmp13354 + r_run_k_29);
	assign w_sys_tmp13354 = 32'sh00001e61;
	assign w_sys_tmp13358 = (w_sys_tmp13359 + r_run_k_29);
	assign w_sys_tmp13359 = 32'sh00001ec6;
	assign w_sys_tmp13363 = (w_sys_tmp13364 + r_run_k_29);
	assign w_sys_tmp13364 = 32'sh00001f2b;
	assign w_sys_tmp13368 = (w_sys_tmp13369 + r_run_k_29);
	assign w_sys_tmp13369 = 32'sh00001f90;
	assign w_sys_tmp13373 = (w_sys_tmp13374 + r_run_k_29);
	assign w_sys_tmp13374 = 32'sh00001ff5;
	assign w_sys_tmp13378 = (w_sys_tmp13379 + r_run_k_29);
	assign w_sys_tmp13379 = 32'sh0000205a;
	assign w_sys_tmp13383 = (w_sys_tmp13384 + r_run_k_29);
	assign w_sys_tmp13384 = 32'sh000020bf;
	assign w_sys_tmp13388 = (w_sys_tmp13389 + r_run_k_29);
	assign w_sys_tmp13389 = 32'sh00002124;
	assign w_sys_tmp13393 = (w_sys_tmp13394 + r_run_k_29);
	assign w_sys_tmp13394 = 32'sh00002189;
	assign w_sys_tmp13398 = (w_sys_tmp13399 + r_run_k_29);
	assign w_sys_tmp13399 = 32'sh000021ee;
	assign w_sys_tmp13403 = (w_sys_tmp13404 + r_run_k_29);
	assign w_sys_tmp13404 = 32'sh00002253;
	assign w_sys_tmp13408 = (w_sys_tmp13409 + r_run_k_29);
	assign w_sys_tmp13409 = 32'sh000022b8;
	assign w_sys_tmp13413 = (w_sys_tmp13414 + r_run_k_29);
	assign w_sys_tmp13414 = 32'sh0000231d;
	assign w_sys_tmp13418 = (w_sys_tmp13419 + r_run_k_29);
	assign w_sys_tmp13419 = 32'sh00002382;
	assign w_sys_tmp13423 = (w_sys_tmp13424 + r_run_k_29);
	assign w_sys_tmp13424 = 32'sh000023e7;
	assign w_sys_tmp13428 = (w_sys_tmp13429 + r_run_k_29);
	assign w_sys_tmp13429 = 32'sh0000244c;
	assign w_sys_tmp13433 = (w_sys_tmp13434 + r_run_k_29);
	assign w_sys_tmp13434 = 32'sh000024b1;
	assign w_sys_tmp13438 = (w_sys_tmp13439 + r_run_k_29);
	assign w_sys_tmp13439 = 32'sh00002516;
	assign w_sys_tmp13443 = (w_sys_tmp13444 + r_run_k_29);
	assign w_sys_tmp13444 = 32'sh0000257b;
	assign w_sys_tmp13448 = (w_sys_tmp13449 + r_run_k_29);
	assign w_sys_tmp13449 = 32'sh000025e0;
	assign w_sys_tmp13453 = (w_sys_tmp13454 + r_run_k_29);
	assign w_sys_tmp13454 = 32'sh00002645;
	assign w_sys_tmp13458 = (w_sys_tmp13459 + r_run_k_29);
	assign w_sys_tmp13459 = 32'sh000026aa;
	assign w_sys_tmp13463 = (w_sys_tmp13464 + r_run_k_29);
	assign w_sys_tmp13464 = 32'sh0000270f;
	assign w_sys_tmp13468 = (w_sys_tmp13469 + r_run_k_29);
	assign w_sys_tmp13469 = 32'sh00002774;
	assign w_sys_tmp13472 = (r_run_k_29 + w_sys_intOne);


	sub19
		sub19_inst(
			.i_fld_T_0_addr_0 (w_sub19_T_addr),
			.i_fld_T_0_datain_0 (w_sub19_T_datain),
			.o_fld_T_0_dataout_0 (w_sub19_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub19_T_r_w),
			.i_fld_U_2_addr_0 (w_sub19_U_addr),
			.i_fld_U_2_datain_0 (w_sub19_U_datain),
			.o_fld_U_2_dataout_0 (w_sub19_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub19_U_r_w),
			.i_fld_V_1_addr_0 (w_sub19_V_addr),
			.i_fld_V_1_datain_0 (w_sub19_V_datain),
			.o_fld_V_1_dataout_0 (w_sub19_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub19_V_r_w),
			.i_fld_result_3_addr_0 (w_sub19_result_addr),
			.i_fld_result_3_datain_0 (w_sub19_result_datain),
			.o_fld_result_3_dataout_0 (w_sub19_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub19_result_r_w),
			.o_run_busy (w_sub19_run_busy),
			.i_run_req (r_sub19_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub09
		sub09_inst(
			.i_fld_T_0_addr_0 (w_sub09_T_addr),
			.i_fld_T_0_datain_0 (w_sub09_T_datain),
			.o_fld_T_0_dataout_0 (w_sub09_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub09_T_r_w),
			.i_fld_U_2_addr_0 (w_sub09_U_addr),
			.i_fld_U_2_datain_0 (w_sub09_U_datain),
			.o_fld_U_2_dataout_0 (w_sub09_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub09_U_r_w),
			.i_fld_V_1_addr_0 (w_sub09_V_addr),
			.i_fld_V_1_datain_0 (w_sub09_V_datain),
			.o_fld_V_1_dataout_0 (w_sub09_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub09_V_r_w),
			.i_fld_result_3_addr_0 (w_sub09_result_addr),
			.i_fld_result_3_datain_0 (w_sub09_result_datain),
			.o_fld_result_3_dataout_0 (w_sub09_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub09_result_r_w),
			.o_run_busy (w_sub09_run_busy),
			.i_run_req (r_sub09_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub08
		sub08_inst(
			.i_fld_T_0_addr_0 (w_sub08_T_addr),
			.i_fld_T_0_datain_0 (w_sub08_T_datain),
			.o_fld_T_0_dataout_0 (w_sub08_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub08_T_r_w),
			.i_fld_U_2_addr_0 (w_sub08_U_addr),
			.i_fld_U_2_datain_0 (w_sub08_U_datain),
			.o_fld_U_2_dataout_0 (w_sub08_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub08_U_r_w),
			.i_fld_V_1_addr_0 (w_sub08_V_addr),
			.i_fld_V_1_datain_0 (w_sub08_V_datain),
			.o_fld_V_1_dataout_0 (w_sub08_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub08_V_r_w),
			.i_fld_result_3_addr_0 (w_sub08_result_addr),
			.i_fld_result_3_datain_0 (w_sub08_result_datain),
			.o_fld_result_3_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub08_result_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub24
		sub24_inst(
			.i_fld_T_0_addr_0 (w_sub24_T_addr),
			.i_fld_T_0_datain_0 (w_sub24_T_datain),
			.o_fld_T_0_dataout_0 (w_sub24_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub24_T_r_w),
			.i_fld_U_2_addr_0 (w_sub24_U_addr),
			.i_fld_U_2_datain_0 (w_sub24_U_datain),
			.o_fld_U_2_dataout_0 (w_sub24_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub24_U_r_w),
			.i_fld_V_1_addr_0 (w_sub24_V_addr),
			.i_fld_V_1_datain_0 (w_sub24_V_datain),
			.o_fld_V_1_dataout_0 (w_sub24_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub24_V_r_w),
			.i_fld_result_3_addr_0 (w_sub24_result_addr),
			.i_fld_result_3_datain_0 (w_sub24_result_datain),
			.o_fld_result_3_dataout_0 (w_sub24_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub24_result_r_w),
			.o_run_busy (w_sub24_run_busy),
			.i_run_req (r_sub24_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub22
		sub22_inst(
			.i_fld_T_0_addr_0 (w_sub22_T_addr),
			.i_fld_T_0_datain_0 (w_sub22_T_datain),
			.o_fld_T_0_dataout_0 (w_sub22_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub22_T_r_w),
			.i_fld_U_2_addr_0 (w_sub22_U_addr),
			.i_fld_U_2_datain_0 (w_sub22_U_datain),
			.o_fld_U_2_dataout_0 (w_sub22_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub22_U_r_w),
			.i_fld_V_1_addr_0 (w_sub22_V_addr),
			.i_fld_V_1_datain_0 (w_sub22_V_datain),
			.o_fld_V_1_dataout_0 (w_sub22_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub22_V_r_w),
			.i_fld_result_3_addr_0 (w_sub22_result_addr),
			.i_fld_result_3_datain_0 (w_sub22_result_datain),
			.o_fld_result_3_dataout_0 (w_sub22_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub22_result_r_w),
			.o_run_busy (w_sub22_run_busy),
			.i_run_req (r_sub22_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub23
		sub23_inst(
			.i_fld_T_0_addr_0 (w_sub23_T_addr),
			.i_fld_T_0_datain_0 (w_sub23_T_datain),
			.o_fld_T_0_dataout_0 (w_sub23_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub23_T_r_w),
			.i_fld_U_2_addr_0 (w_sub23_U_addr),
			.i_fld_U_2_datain_0 (w_sub23_U_datain),
			.o_fld_U_2_dataout_0 (w_sub23_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub23_U_r_w),
			.i_fld_V_1_addr_0 (w_sub23_V_addr),
			.i_fld_V_1_datain_0 (w_sub23_V_datain),
			.o_fld_V_1_dataout_0 (w_sub23_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub23_V_r_w),
			.i_fld_result_3_addr_0 (w_sub23_result_addr),
			.i_fld_result_3_datain_0 (w_sub23_result_datain),
			.o_fld_result_3_dataout_0 (w_sub23_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub23_result_r_w),
			.o_run_busy (w_sub23_run_busy),
			.i_run_req (r_sub23_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub12
		sub12_inst(
			.i_fld_T_0_addr_0 (w_sub12_T_addr),
			.i_fld_T_0_datain_0 (w_sub12_T_datain),
			.o_fld_T_0_dataout_0 (w_sub12_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub12_T_r_w),
			.i_fld_U_2_addr_0 (w_sub12_U_addr),
			.i_fld_U_2_datain_0 (w_sub12_U_datain),
			.o_fld_U_2_dataout_0 (w_sub12_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub12_U_r_w),
			.i_fld_V_1_addr_0 (w_sub12_V_addr),
			.i_fld_V_1_datain_0 (w_sub12_V_datain),
			.o_fld_V_1_dataout_0 (w_sub12_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub12_V_r_w),
			.i_fld_result_3_addr_0 (w_sub12_result_addr),
			.i_fld_result_3_datain_0 (w_sub12_result_datain),
			.o_fld_result_3_dataout_0 (w_sub12_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub12_result_r_w),
			.o_run_busy (w_sub12_run_busy),
			.i_run_req (r_sub12_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_T_0_addr_0 (w_sub03_T_addr),
			.i_fld_T_0_datain_0 (w_sub03_T_datain),
			.o_fld_T_0_dataout_0 (w_sub03_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub03_T_r_w),
			.i_fld_U_2_addr_0 (w_sub03_U_addr),
			.i_fld_U_2_datain_0 (w_sub03_U_datain),
			.o_fld_U_2_dataout_0 (w_sub03_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub03_U_r_w),
			.i_fld_V_1_addr_0 (w_sub03_V_addr),
			.i_fld_V_1_datain_0 (w_sub03_V_datain),
			.o_fld_V_1_dataout_0 (w_sub03_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub03_V_r_w),
			.i_fld_result_3_addr_0 (w_sub03_result_addr),
			.i_fld_result_3_datain_0 (w_sub03_result_datain),
			.o_fld_result_3_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub03_result_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_T_0_addr_0 (w_sub02_T_addr),
			.i_fld_T_0_datain_0 (w_sub02_T_datain),
			.o_fld_T_0_dataout_0 (w_sub02_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub02_T_r_w),
			.i_fld_U_2_addr_0 (w_sub02_U_addr),
			.i_fld_U_2_datain_0 (w_sub02_U_datain),
			.o_fld_U_2_dataout_0 (w_sub02_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub02_U_r_w),
			.i_fld_V_1_addr_0 (w_sub02_V_addr),
			.i_fld_V_1_datain_0 (w_sub02_V_datain),
			.o_fld_V_1_dataout_0 (w_sub02_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub02_V_r_w),
			.i_fld_result_3_addr_0 (w_sub02_result_addr),
			.i_fld_result_3_datain_0 (w_sub02_result_datain),
			.o_fld_result_3_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub02_result_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub11
		sub11_inst(
			.i_fld_T_0_addr_0 (w_sub11_T_addr),
			.i_fld_T_0_datain_0 (w_sub11_T_datain),
			.o_fld_T_0_dataout_0 (w_sub11_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub11_T_r_w),
			.i_fld_U_2_addr_0 (w_sub11_U_addr),
			.i_fld_U_2_datain_0 (w_sub11_U_datain),
			.o_fld_U_2_dataout_0 (w_sub11_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub11_U_r_w),
			.i_fld_V_1_addr_0 (w_sub11_V_addr),
			.i_fld_V_1_datain_0 (w_sub11_V_datain),
			.o_fld_V_1_dataout_0 (w_sub11_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub11_V_r_w),
			.i_fld_result_3_addr_0 (w_sub11_result_addr),
			.i_fld_result_3_datain_0 (w_sub11_result_datain),
			.o_fld_result_3_dataout_0 (w_sub11_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub11_result_r_w),
			.o_run_busy (w_sub11_run_busy),
			.i_run_req (r_sub11_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub14
		sub14_inst(
			.i_fld_T_0_addr_0 (w_sub14_T_addr),
			.i_fld_T_0_datain_0 (w_sub14_T_datain),
			.o_fld_T_0_dataout_0 (w_sub14_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub14_T_r_w),
			.i_fld_U_2_addr_0 (w_sub14_U_addr),
			.i_fld_U_2_datain_0 (w_sub14_U_datain),
			.o_fld_U_2_dataout_0 (w_sub14_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub14_U_r_w),
			.i_fld_V_1_addr_0 (w_sub14_V_addr),
			.i_fld_V_1_datain_0 (w_sub14_V_datain),
			.o_fld_V_1_dataout_0 (w_sub14_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub14_V_r_w),
			.i_fld_result_3_addr_0 (w_sub14_result_addr),
			.i_fld_result_3_datain_0 (w_sub14_result_datain),
			.o_fld_result_3_dataout_0 (w_sub14_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub14_result_r_w),
			.o_run_busy (w_sub14_run_busy),
			.i_run_req (r_sub14_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_T_0_addr_0 (w_sub01_T_addr),
			.i_fld_T_0_datain_0 (w_sub01_T_datain),
			.o_fld_T_0_dataout_0 (w_sub01_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub01_T_r_w),
			.i_fld_U_2_addr_0 (w_sub01_U_addr),
			.i_fld_U_2_datain_0 (w_sub01_U_datain),
			.o_fld_U_2_dataout_0 (w_sub01_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub01_U_r_w),
			.i_fld_V_1_addr_0 (w_sub01_V_addr),
			.i_fld_V_1_datain_0 (w_sub01_V_datain),
			.o_fld_V_1_dataout_0 (w_sub01_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub01_V_r_w),
			.i_fld_result_3_addr_0 (w_sub01_result_addr),
			.i_fld_result_3_datain_0 (w_sub01_result_datain),
			.o_fld_result_3_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub01_result_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_T_0_addr_0 (w_sub00_T_addr),
			.i_fld_T_0_datain_0 (w_sub00_T_datain),
			.o_fld_T_0_dataout_0 (w_sub00_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub00_T_r_w),
			.i_fld_U_2_addr_0 (w_sub00_U_addr),
			.i_fld_U_2_datain_0 (w_sub00_U_datain),
			.o_fld_U_2_dataout_0 (w_sub00_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub00_U_r_w),
			.i_fld_V_1_addr_0 (w_sub00_V_addr),
			.i_fld_V_1_datain_0 (w_sub00_V_datain),
			.o_fld_V_1_dataout_0 (w_sub00_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub00_V_r_w),
			.i_fld_result_3_addr_0 (w_sub00_result_addr),
			.i_fld_result_3_datain_0 (w_sub00_result_datain),
			.o_fld_result_3_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub00_result_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub13
		sub13_inst(
			.i_fld_T_0_addr_0 (w_sub13_T_addr),
			.i_fld_T_0_datain_0 (w_sub13_T_datain),
			.o_fld_T_0_dataout_0 (w_sub13_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub13_T_r_w),
			.i_fld_U_2_addr_0 (w_sub13_U_addr),
			.i_fld_U_2_datain_0 (w_sub13_U_datain),
			.o_fld_U_2_dataout_0 (w_sub13_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub13_U_r_w),
			.i_fld_V_1_addr_0 (w_sub13_V_addr),
			.i_fld_V_1_datain_0 (w_sub13_V_datain),
			.o_fld_V_1_dataout_0 (w_sub13_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub13_V_r_w),
			.i_fld_result_3_addr_0 (w_sub13_result_addr),
			.i_fld_result_3_datain_0 (w_sub13_result_datain),
			.o_fld_result_3_dataout_0 (w_sub13_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub13_result_r_w),
			.o_run_busy (w_sub13_run_busy),
			.i_run_req (r_sub13_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_T_0_addr_0 (w_sub07_T_addr),
			.i_fld_T_0_datain_0 (w_sub07_T_datain),
			.o_fld_T_0_dataout_0 (w_sub07_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub07_T_r_w),
			.i_fld_U_2_addr_0 (w_sub07_U_addr),
			.i_fld_U_2_datain_0 (w_sub07_U_datain),
			.o_fld_U_2_dataout_0 (w_sub07_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub07_U_r_w),
			.i_fld_V_1_addr_0 (w_sub07_V_addr),
			.i_fld_V_1_datain_0 (w_sub07_V_datain),
			.o_fld_V_1_dataout_0 (w_sub07_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub07_V_r_w),
			.i_fld_result_3_addr_0 (w_sub07_result_addr),
			.i_fld_result_3_datain_0 (w_sub07_result_datain),
			.o_fld_result_3_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub07_result_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub16
		sub16_inst(
			.i_fld_T_0_addr_0 (w_sub16_T_addr),
			.i_fld_T_0_datain_0 (w_sub16_T_datain),
			.o_fld_T_0_dataout_0 (w_sub16_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub16_T_r_w),
			.i_fld_U_2_addr_0 (w_sub16_U_addr),
			.i_fld_U_2_datain_0 (w_sub16_U_datain),
			.o_fld_U_2_dataout_0 (w_sub16_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub16_U_r_w),
			.i_fld_V_1_addr_0 (w_sub16_V_addr),
			.i_fld_V_1_datain_0 (w_sub16_V_datain),
			.o_fld_V_1_dataout_0 (w_sub16_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub16_V_r_w),
			.i_fld_result_3_addr_0 (w_sub16_result_addr),
			.i_fld_result_3_datain_0 (w_sub16_result_datain),
			.o_fld_result_3_dataout_0 (w_sub16_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub16_result_r_w),
			.o_run_busy (w_sub16_run_busy),
			.i_run_req (r_sub16_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_T_0_addr_0 (w_sub06_T_addr),
			.i_fld_T_0_datain_0 (w_sub06_T_datain),
			.o_fld_T_0_dataout_0 (w_sub06_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub06_T_r_w),
			.i_fld_U_2_addr_0 (w_sub06_U_addr),
			.i_fld_U_2_datain_0 (w_sub06_U_datain),
			.o_fld_U_2_dataout_0 (w_sub06_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub06_U_r_w),
			.i_fld_V_1_addr_0 (w_sub06_V_addr),
			.i_fld_V_1_datain_0 (w_sub06_V_datain),
			.o_fld_V_1_dataout_0 (w_sub06_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub06_V_r_w),
			.i_fld_result_3_addr_0 (w_sub06_result_addr),
			.i_fld_result_3_datain_0 (w_sub06_result_datain),
			.o_fld_result_3_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub06_result_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub15
		sub15_inst(
			.i_fld_T_0_addr_0 (w_sub15_T_addr),
			.i_fld_T_0_datain_0 (w_sub15_T_datain),
			.o_fld_T_0_dataout_0 (w_sub15_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub15_T_r_w),
			.i_fld_U_2_addr_0 (w_sub15_U_addr),
			.i_fld_U_2_datain_0 (w_sub15_U_datain),
			.o_fld_U_2_dataout_0 (w_sub15_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub15_U_r_w),
			.i_fld_V_1_addr_0 (w_sub15_V_addr),
			.i_fld_V_1_datain_0 (w_sub15_V_datain),
			.o_fld_V_1_dataout_0 (w_sub15_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub15_V_r_w),
			.i_fld_result_3_addr_0 (w_sub15_result_addr),
			.i_fld_result_3_datain_0 (w_sub15_result_datain),
			.o_fld_result_3_dataout_0 (w_sub15_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub15_result_r_w),
			.o_run_busy (w_sub15_run_busy),
			.i_run_req (r_sub15_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_T_0_addr_0 (w_sub05_T_addr),
			.i_fld_T_0_datain_0 (w_sub05_T_datain),
			.o_fld_T_0_dataout_0 (w_sub05_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub05_T_r_w),
			.i_fld_U_2_addr_0 (w_sub05_U_addr),
			.i_fld_U_2_datain_0 (w_sub05_U_datain),
			.o_fld_U_2_dataout_0 (w_sub05_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub05_U_r_w),
			.i_fld_V_1_addr_0 (w_sub05_V_addr),
			.i_fld_V_1_datain_0 (w_sub05_V_datain),
			.o_fld_V_1_dataout_0 (w_sub05_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub05_V_r_w),
			.i_fld_result_3_addr_0 (w_sub05_result_addr),
			.i_fld_result_3_datain_0 (w_sub05_result_datain),
			.o_fld_result_3_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub05_result_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub18
		sub18_inst(
			.i_fld_T_0_addr_0 (w_sub18_T_addr),
			.i_fld_T_0_datain_0 (w_sub18_T_datain),
			.o_fld_T_0_dataout_0 (w_sub18_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub18_T_r_w),
			.i_fld_U_2_addr_0 (w_sub18_U_addr),
			.i_fld_U_2_datain_0 (w_sub18_U_datain),
			.o_fld_U_2_dataout_0 (w_sub18_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub18_U_r_w),
			.i_fld_V_1_addr_0 (w_sub18_V_addr),
			.i_fld_V_1_datain_0 (w_sub18_V_datain),
			.o_fld_V_1_dataout_0 (w_sub18_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub18_V_r_w),
			.i_fld_result_3_addr_0 (w_sub18_result_addr),
			.i_fld_result_3_datain_0 (w_sub18_result_datain),
			.o_fld_result_3_dataout_0 (w_sub18_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub18_result_r_w),
			.o_run_busy (w_sub18_run_busy),
			.i_run_req (r_sub18_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_T_0_addr_0 (w_sub04_T_addr),
			.i_fld_T_0_datain_0 (w_sub04_T_datain),
			.o_fld_T_0_dataout_0 (w_sub04_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub04_T_r_w),
			.i_fld_U_2_addr_0 (w_sub04_U_addr),
			.i_fld_U_2_datain_0 (w_sub04_U_datain),
			.o_fld_U_2_dataout_0 (w_sub04_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub04_U_r_w),
			.i_fld_V_1_addr_0 (w_sub04_V_addr),
			.i_fld_V_1_datain_0 (w_sub04_V_datain),
			.o_fld_V_1_dataout_0 (w_sub04_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub04_V_r_w),
			.i_fld_result_3_addr_0 (w_sub04_result_addr),
			.i_fld_result_3_datain_0 (w_sub04_result_datain),
			.o_fld_result_3_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub04_result_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub17
		sub17_inst(
			.i_fld_T_0_addr_0 (w_sub17_T_addr),
			.i_fld_T_0_datain_0 (w_sub17_T_datain),
			.o_fld_T_0_dataout_0 (w_sub17_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub17_T_r_w),
			.i_fld_U_2_addr_0 (w_sub17_U_addr),
			.i_fld_U_2_datain_0 (w_sub17_U_datain),
			.o_fld_U_2_dataout_0 (w_sub17_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub17_U_r_w),
			.i_fld_V_1_addr_0 (w_sub17_V_addr),
			.i_fld_V_1_datain_0 (w_sub17_V_datain),
			.o_fld_V_1_dataout_0 (w_sub17_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub17_V_r_w),
			.i_fld_result_3_addr_0 (w_sub17_result_addr),
			.i_fld_result_3_datain_0 (w_sub17_result_datain),
			.o_fld_result_3_dataout_0 (w_sub17_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub17_result_r_w),
			.o_run_busy (w_sub17_run_busy),
			.i_run_req (r_sub17_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub10
		sub10_inst(
			.i_fld_T_0_addr_0 (w_sub10_T_addr),
			.i_fld_T_0_datain_0 (w_sub10_T_datain),
			.o_fld_T_0_dataout_0 (w_sub10_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub10_T_r_w),
			.i_fld_U_2_addr_0 (w_sub10_U_addr),
			.i_fld_U_2_datain_0 (w_sub10_U_datain),
			.o_fld_U_2_dataout_0 (w_sub10_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub10_U_r_w),
			.i_fld_V_1_addr_0 (w_sub10_V_addr),
			.i_fld_V_1_datain_0 (w_sub10_V_datain),
			.o_fld_V_1_dataout_0 (w_sub10_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub10_V_r_w),
			.i_fld_result_3_addr_0 (w_sub10_result_addr),
			.i_fld_result_3_datain_0 (w_sub10_result_datain),
			.o_fld_result_3_dataout_0 (w_sub10_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub10_result_r_w),
			.o_run_busy (w_sub10_run_busy),
			.i_run_req (r_sub10_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub20
		sub20_inst(
			.i_fld_T_0_addr_0 (w_sub20_T_addr),
			.i_fld_T_0_datain_0 (w_sub20_T_datain),
			.o_fld_T_0_dataout_0 (w_sub20_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub20_T_r_w),
			.i_fld_U_2_addr_0 (w_sub20_U_addr),
			.i_fld_U_2_datain_0 (w_sub20_U_datain),
			.o_fld_U_2_dataout_0 (w_sub20_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub20_U_r_w),
			.i_fld_V_1_addr_0 (w_sub20_V_addr),
			.i_fld_V_1_datain_0 (w_sub20_V_datain),
			.o_fld_V_1_dataout_0 (w_sub20_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub20_V_r_w),
			.i_fld_result_3_addr_0 (w_sub20_result_addr),
			.i_fld_result_3_datain_0 (w_sub20_result_datain),
			.o_fld_result_3_dataout_0 (w_sub20_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub20_result_r_w),
			.o_run_busy (w_sub20_run_busy),
			.i_run_req (r_sub20_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub21
		sub21_inst(
			.i_fld_T_0_addr_0 (w_sub21_T_addr),
			.i_fld_T_0_datain_0 (w_sub21_T_datain),
			.o_fld_T_0_dataout_0 (w_sub21_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub21_T_r_w),
			.i_fld_U_2_addr_0 (w_sub21_U_addr),
			.i_fld_U_2_datain_0 (w_sub21_U_datain),
			.o_fld_U_2_dataout_0 (w_sub21_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub21_U_r_w),
			.i_fld_V_1_addr_0 (w_sub21_V_addr),
			.i_fld_V_1_datain_0 (w_sub21_V_datain),
			.o_fld_V_1_dataout_0 (w_sub21_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub21_V_r_w),
			.i_fld_result_3_addr_0 (w_sub21_result_addr),
			.i_fld_result_3_datain_0 (w_sub21_result_datain),
			.o_fld_result_3_dataout_0 (w_sub21_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub21_result_r_w),
			.o_run_busy (w_sub21_run_busy),
			.i_run_req (r_sub21_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(14), .WORDS(10404) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(14), .WORDS(10404) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(14), .WORDS(10404) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(14), .WORDS(10404) )
		dpram_V_3(
			.clk (clock),
			.ce_0 (w_fld_V_3_ce_0),
			.addr_0 (w_fld_V_3_addr_0),
			.datain_0 (w_fld_V_3_datain_0),
			.dataout_0 (w_fld_V_3_dataout_0),
			.r_w_0 (w_fld_V_3_r_w_0),
			.ce_1 (w_fld_V_3_ce_1),
			.addr_1 (r_fld_V_3_addr_1),
			.datain_1 (r_fld_V_3_datain_1),
			.dataout_1 (w_fld_V_3_dataout_1),
			.r_w_1 (r_fld_V_3_r_w_1)
		);

	DivInt
		DivInt_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.dividend (r_ip_DivInt_dividend_0),
			.divisor (r_ip_DivInt_divisor_0),
			.fractional (w_ip_DivInt_fractional_0),
			.quotient (w_ip_DivInt_quotient_0)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_ip_DivInt_dividend_0 <= r_run_mx_32;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_ip_DivInt_dividend_0 <= r_run_mx_32;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_ip_DivInt_divisor_0 <= w_sys_tmp7319;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_ip_DivInt_divisor_0 <= w_sys_tmp7323;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h27) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h33) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h3b)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp38;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h33)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp297[31], w_sys_tmp297[30:0] };

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp269[31], w_sys_tmp269[30:0] };

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp297[31], w_sys_tmp297[30:0] };

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp269[31], w_sys_tmp269[30:0] };

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp185[31], w_sys_tmp185[30:0] };

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp185[31], w_sys_tmp185[30:0] };

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp269[31], w_sys_tmp269[30:0] };

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp297[31], w_sys_tmp297[30:0] };

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp269[31], w_sys_tmp269[30:0] };

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp297[31], w_sys_tmp297[30:0] };

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp157[31], w_sys_tmp157[30:0] };

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp185[31], w_sys_tmp185[30:0] };

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp185[31], w_sys_tmp185[30:0] };

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp128[31], w_sys_tmp128[30:0] };

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp213[31], w_sys_tmp213[30:0] };

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp37[31], w_sys_tmp37[30:0] };

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp185[31], w_sys_tmp185[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h2f) || (r_sys_run_step==9'h36) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h41)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==9'hc) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h27) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h33) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h3d)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp36;

									end
									else
									if((r_sys_run_step==9'h20) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h32) || (r_sys_run_step==9'h38)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==9'h1a) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h3e) || (r_sys_run_step==9'h40)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp16_float;

									end
									else
									if((9'h7<=r_sys_run_step && r_sys_run_step<=9'hb) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h31)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_36;

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h1f)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==9'hd) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h2e)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==9'h17) || (r_sys_run_step==9'h28)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp37;

									end
									else
									if((r_sys_run_step==9'h1a) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h32) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h42)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==9'h23) || (r_sys_run_step==9'h2f) || (r_sys_run_step==9'h38)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==9'h16) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h36) || (r_sys_run_step==9'h3e) || (r_sys_run_step==9'h41)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==9'he) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h27) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h33) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h3d)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_41;

									end
									else
									if((9'h7<=r_sys_run_step && r_sys_run_step<=9'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==9'h1d) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h3c) || (r_sys_run_step==9'h40)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp11_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp20;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp15) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h47)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp588) ? 7'h13 : 7'h15);

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1af)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp5754) ? 7'h19 : 7'h1b);

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6d)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7055) ? 7'h20 : 7'h4d);

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7058) ? 7'h24 : 7'h26);

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7075) ? 7'h2a : 7'h2c);

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h27)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h25)) begin
										r_sys_run_phase <= ((w_sys_tmp7320) ? 7'h30 : 7'h32);

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp7445) ? 7'h36 : 7'h38);

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b5)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10067) ? 7'h3c : 7'h3d);

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6e)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_phase <= 7'h3f;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_phase <= 7'h41;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h42;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp10727) ? 7'h45 : 7'h47);

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b9)) begin
										r_sys_run_phase <= 7'h42;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= 7'h48;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp12953) ? 7'h4b : 7'h1d);

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h64)) begin
										r_sys_run_phase <= 7'h48;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 5'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h47)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1af)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6d)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h27)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h25)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h25)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b5)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6e)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b9)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h64)) begin
										r_sys_run_stage <= 5'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 9'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h47)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h46)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1af)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1ae)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6d)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6c)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h1) || (r_sys_run_step==9'h2)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h27)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h26)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h25)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h25)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h24)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h12)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b5)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1b4)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6e)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6d)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub09_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub10_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub11_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub12_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub13_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub14_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub15_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub16_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub17_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub18_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub19_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub20_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub21_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub22_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub23_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h1)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= ((w_sub24_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1b8)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==9'h1b9)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sys_run_step <= 9'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h64)) begin
										r_sys_run_step <= 9'h0;

									end
									else
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h63)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h4d: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp22[13:0] );

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7066[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7070[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7062[13:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h2) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7079[13:0] );

									end
									else
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h3) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7084[13:0] );

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7326[13:0] );

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7690[13:0] );

									end
									else
									if((r_sys_run_step==9'h14) || (r_sys_run_step==9'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7570[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7642[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8104[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ab)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10012[13:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8794[13:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9316[13:0] );

									end
									else
									if((r_sys_run_step==9'h98) || (r_sys_run_step==9'h9a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8362[13:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9694[13:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8350[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9988[13:0] );

									end
									else
									if((r_sys_run_step==9'h197)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9892[13:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8524[13:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8578[13:0] );

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9478[13:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9622[13:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8122[13:0] );

									end
									else
									if((r_sys_run_step==9'h182)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9766[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7810[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9976[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7750[13:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9052[13:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8602[13:0] );

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8998[13:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9334[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7504[13:0] );

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9640[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10048[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7672[13:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9058[13:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9202[13:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8458[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7486[13:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9736[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8044[13:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9454[13:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8380[13:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8284[13:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8548[13:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8908[13:0] );

									end
									else
									if((r_sys_run_step==9'h192)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9862[13:0] );

									end
									else
									if((r_sys_run_step==9'h40) || (r_sys_run_step==9'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7834[13:0] );

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9340[13:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9118[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7492[13:0] );

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8866[13:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8926[13:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8836[13:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9442[13:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8554[13:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8182[13:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9526[13:0] );

									end
									else
									if((r_sys_run_step==9'h171) || (r_sys_run_step==9'h173)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9664[13:0] );

									end
									else
									if((r_sys_run_step==9'h187) || (r_sys_run_step==9'h189)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9796[13:0] );

									end
									else
									if((r_sys_run_step==9'h19b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9916[13:0] );

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8872[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7702[13:0] );

									end
									else
									if((r_sys_run_step==9'h41) || (r_sys_run_step==9'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7840[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7990[13:0] );

									end
									else
									if((r_sys_run_step==9'h130) || (r_sys_run_step==9'h132)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9274[13:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8422[13:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9358[13:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8800[13:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8962[13:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9838[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9970[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ae)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10030[13:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8326[13:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9382[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7822[13:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9100[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7450[13:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9658[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7516[13:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8272[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8026[13:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9406[13:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8410[13:0] );

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9568[13:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8314[13:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9106[13:0] );

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8446[13:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8398[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8002[13:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9514[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7948[13:0] );

									end
									else
									if((r_sys_run_step==9'h104) || (r_sys_run_step==9'h106)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9010[13:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8752[13:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8608[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7828[13:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8644[13:0] );

									end
									else
									if((r_sys_run_step==9'h82) || (r_sys_run_step==9'h84)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8230[13:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8788[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7762[13:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8764[13:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9730[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7732[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7918[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7522[13:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8170[13:0] );

									end
									else
									if((r_sys_run_step==9'h12d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9256[13:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8596[13:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8206[13:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9298[13:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8296[13:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9064[13:0] );

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9856[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7738[13:0] );

									end
									else
									if((r_sys_run_step==9'hee) || (r_sys_run_step==9'hf0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8878[13:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9034[13:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9046[13:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8164[13:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9574[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ad)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10024[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9964[13:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9310[13:0] );

									end
									else
									if((r_sys_run_step==9'h15c) || (r_sys_run_step==9'h15e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9538[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7882[13:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8848[13:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9586[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7912[13:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9364[13:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8824[13:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8260[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7942[13:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9436[13:0] );

									end
									else
									if((r_sys_run_step==9'h199)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9904[13:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8914[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7924[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7906[13:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8110[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7888[13:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8842[13:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8464[13:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8152[13:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9448[13:0] );

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9124[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7900[13:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8308[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9994[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7534[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7600[13:0] );

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9244[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8092[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10060[13:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8482[13:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9322[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7798[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7606[13:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9868[13:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8140[13:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9226[13:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8470[13:0] );

									end
									else
									if((r_sys_run_step==9'hae) || (r_sys_run_step==9'hb0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8494[13:0] );

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8668[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ac)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10018[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7960[13:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9424[13:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8434[13:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8950[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7540[13:0] );

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9502[13:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8176[13:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8212[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7756[13:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8542[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7678[13:0] );

									end
									else
									if((r_sys_run_step==9'h131) || (r_sys_run_step==9'h133)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9280[13:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8704[13:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8566[13:0] );

									end
									else
									if((r_sys_run_step==9'h188) || (r_sys_run_step==9'h18a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9802[13:0] );

									end
									else
									if((r_sys_run_step==9'h157)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9508[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7876[13:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9040[13:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8686[13:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8734[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7618[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7696[13:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9214[13:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8254[13:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8944[13:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8920[13:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8698[13:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8932[13:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9094[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8062[13:0] );

									end
									else
									if((r_sys_run_step==9'h81) || (r_sys_run_step==9'h83)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8224[13:0] );

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9460[13:0] );

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8854[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8080[13:0] );

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9466[13:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8098[13:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8902[13:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8776[13:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8158[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8086[13:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9724[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7594[13:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8512[13:0] );

									end
									else
									if((r_sys_run_step==9'h15) || (r_sys_run_step==9'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7576[13:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9370[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7996[13:0] );

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9646[13:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9208[13:0] );

									end
									else
									if((r_sys_run_step==9'h1af)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10036[13:0] );

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9130[13:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9712[13:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8716[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7894[13:0] );

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8986[13:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8218[13:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9394[13:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9352[13:0] );

									end
									else
									if((r_sys_run_step==9'h11a) || (r_sys_run_step==9'h11c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9142[13:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9718[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10000[13:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8830[13:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9556[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7666[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7612[13:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9328[13:0] );

									end
									else
									if((r_sys_run_step==9'h19c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9922[13:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8248[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8074[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7660[13:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8290[13:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8404[13:0] );

									end
									else
									if((r_sys_run_step==9'hc4) || (r_sys_run_step==9'hc6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8626[13:0] );

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9250[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7744[13:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8116[13:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8440[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7624[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7774[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8008[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7654[13:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8338[13:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8134[13:0] );

									end
									else
									if((r_sys_run_step==9'h1aa)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10006[13:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8536[13:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9592[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8050[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7792[13:0] );

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9634[13:0] );

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9472[13:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8572[13:0] );

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8656[13:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9820[13:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9196[13:0] );

									end
									else
									if((r_sys_run_step==9'h15b) || (r_sys_run_step==9'h15d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9532[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7510[13:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9184[13:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9580[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7528[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7708[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7558[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7648[13:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9616[13:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9088[13:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9562[13:0] );

									end
									else
									if((r_sys_run_step==9'h97) || (r_sys_run_step==9'h99)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8356[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7954[13:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8320[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7786[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8014[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7864[13:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9706[13:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9178[13:0] );

									end
									else
									if((r_sys_run_step==9'h183)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9772[13:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9232[13:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9784[13:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9190[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7636[13:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9844[13:0] );

									end
									else
									if((r_sys_run_step==9'h172) || (r_sys_run_step==9'h174)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9670[13:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8332[13:0] );

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8662[13:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8650[13:0] );

									end
									else
									if((r_sys_run_step==9'hc3) || (r_sys_run_step==9'hc5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8620[13:0] );

									end
									else
									if((r_sys_run_step==9'h19e) || (r_sys_run_step==9'h1a0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9934[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7684[13:0] );

									end
									else
									if((r_sys_run_step==9'h56) || (r_sys_run_step==9'h58)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7966[13:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9376[13:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9790[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7816[13:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9754[13:0] );

									end
									else
									if((r_sys_run_step==9'h19a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9910[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7930[13:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8758[13:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8476[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7780[13:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9430[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7564[13:0] );

									end
									else
									if((r_sys_run_step==9'hef) || (r_sys_run_step==9'hf1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8884[13:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9136[13:0] );

									end
									else
									if((r_sys_run_step==9'had) || (r_sys_run_step==9'haf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8488[13:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8968[13:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8302[13:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9346[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9982[13:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9418[13:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8728[13:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8584[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7468[13:0] );

									end
									else
									if((r_sys_run_step==9'h105) || (r_sys_run_step==9'h107)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9016[13:0] );

									end
									else
									if((r_sys_run_step==9'h12e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9262[13:0] );

									end
									else
									if((r_sys_run_step==9'h57) || (r_sys_run_step==9'h59)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7972[13:0] );

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9004[13:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9220[13:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9700[13:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9166[13:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8722[13:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8770[13:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9688[13:0] );

									end
									else
									if((r_sys_run_step==9'h181)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9760[13:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9400[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8032[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7456[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7858[13:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8146[13:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8974[13:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9238[13:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9604[13:0] );

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8614[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7726[13:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8710[13:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8680[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9958[13:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9832[13:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8590[13:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9070[13:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9112[13:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9652[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10054[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9952[13:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8746[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7462[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7804[13:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8518[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7546[13:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8740[13:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9826[13:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8806[13:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8266[13:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8674[13:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9388[13:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8392[13:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8818[13:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9742[13:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8128[13:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9598[13:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8938[13:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8992[13:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8386[13:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8956[13:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8194[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7936[13:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9610[13:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8980[13:0] );

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9268[13:0] );

									end
									else
									if((r_sys_run_step==9'h195)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9880[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7870[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8056[13:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8812[13:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9412[13:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9172[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8020[13:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8428[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8038[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8068[13:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9748[13:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8782[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7630[13:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8188[13:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8344[13:0] );

									end
									else
									if((r_sys_run_step==9'h11b) || (r_sys_run_step==9'h11d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9148[13:0] );

									end
									else
									if((r_sys_run_step==9'h19d) || (r_sys_run_step==9'h19f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9928[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7768[13:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8452[13:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9496[13:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9850[13:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8530[13:0] );

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9628[13:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8278[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7474[13:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8692[13:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8560[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7498[13:0] );

									end
									else
									if((r_sys_run_step==9'heb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8860[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10042[13:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9076[13:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9484[13:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9490[13:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9520[13:0] );

									end
									else
									if((r_sys_run_step==9'h198)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9898[13:0] );

									end
									else
									if((r_sys_run_step==9'h184)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9778[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7552[13:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9304[13:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8200[13:0] );

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9874[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp7480[13:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp8416[13:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9082[13:0] );

									end
									else
									if((r_sys_run_step==9'h196)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp9886[13:0] );

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10642[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10258[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10522[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10384[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10126[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10660[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10576[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10498[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10552[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10180[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10444[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10408[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10234[13:0] );

									end
									else
									if((r_sys_run_step==9'h14) || (r_sys_run_step==9'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10192[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10270[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10648[13:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10720[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10492[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10540[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10132[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10360[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10516[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10612[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10618[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10450[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10318[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10240[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10558[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10528[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10264[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10324[13:0] );

									end
									else
									if((r_sys_run_step==9'h57) || (r_sys_run_step==9'h59)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10594[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10672[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10216[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10654[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10330[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10348[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10156[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10144[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10570[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10300[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10510[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10684[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10582[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10666[13:0] );

									end
									else
									if((r_sys_run_step==9'h40) || (r_sys_run_step==9'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10456[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10546[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10186[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10102[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10072[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10534[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10168[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10120[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10150[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10390[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10078[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10378[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10276[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10246[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10564[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10114[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10090[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10624[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10438[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10138[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10690[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10228[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10396[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10486[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10084[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10306[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10402[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10678[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10702[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10696[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10366[13:0] );

									end
									else
									if((r_sys_run_step==9'h15) || (r_sys_run_step==9'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10198[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10096[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10222[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10288[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10294[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10630[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10480[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10708[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10108[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10354[13:0] );

									end
									else
									if((r_sys_run_step==9'h56) || (r_sys_run_step==9'h58)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10588[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10426[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10312[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10504[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10162[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10372[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10414[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10252[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10174[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10282[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10714[13:0] );

									end
									else
									if((r_sys_run_step==9'h41) || (r_sys_run_step==9'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10462[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10432[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10636[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10420[13:0] );

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11522[13:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11652[13:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11302[13:0] );

									end
									else
									if((r_sys_run_step==9'h197)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12777[13:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11282[13:0] );

									end
									else
									if((r_sys_run_step==9'h7c) || (r_sys_run_step==9'h7d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11362[13:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12617[13:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11177[13:0] );

									end
									else
									if((r_sys_run_step==9'h26) || (r_sys_run_step==9'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10932[13:0] );

									end
									else
									if((r_sys_run_step==9'h27) || (r_sys_run_step==9'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10937[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11267[13:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11417[13:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11887[13:0] );

									end
									else
									if((r_sys_run_step==9'hc) || (r_sys_run_step==9'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10792[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11232[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11287[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12942[13:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11702[13:0] );

									end
									else
									if((r_sys_run_step==9'h29) || (r_sys_run_step==9'h45)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10947[13:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12537[13:0] );

									end
									else
									if((r_sys_run_step==9'h198)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12782[13:0] );

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12152[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11272[13:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12307[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ae)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12892[13:0] );

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12567[13:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11762[13:0] );

									end
									else
									if((r_sys_run_step==9'h14) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h3e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10840[13:0] );

									end
									else
									if((r_sys_run_step==9'h1aa)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12872[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12937[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12927[13:0] );

									end
									else
									if((r_sys_run_step==9'h15) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10846[13:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11477[13:0] );

									end
									else
									if((r_sys_run_step==9'hd) || (r_sys_run_step==9'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10798[13:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11547[13:0] );

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11502[13:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12382[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11207[13:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11512[13:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12447[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12862[13:0] );

									end
									else
									if((r_sys_run_step==9'h188)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12702[13:0] );

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11757[13:0] );

									end
									else
									if((r_sys_run_step==9'h13) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h3d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10834[13:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12277[13:0] );

									end
									else
									if((r_sys_run_step==9'h196)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12772[13:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11317[13:0] );

									end
									else
									if((r_sys_run_step==9'h19b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12797[13:0] );

									end
									else
									if((r_sys_run_step==9'h19f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12817[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10732[13:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12442[13:0] );

									end
									else
									if((r_sys_run_step==9'h195)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12767[13:0] );

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11927[13:0] );

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12022[13:0] );

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12747[13:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11622[13:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11422[13:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12027[13:0] );

									end
									else
									if((r_sys_run_step==9'h12) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10828[13:0] );

									end
									else
									if((r_sys_run_step==9'h19d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12807[13:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11327[13:0] );

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12562[13:0] );

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11572[13:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11777[13:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12157[13:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12462[13:0] );

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12162[13:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11867[13:0] );

									end
									else
									if((r_sys_run_step==9'h28) || (r_sys_run_step==9'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10942[13:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11877[13:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11582[13:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11432[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12822[13:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11992[13:0] );

									end
									else
									if((r_sys_run_step==9'h32) || (r_sys_run_step==9'h4e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10992[13:0] );

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12427[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10738[13:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12652[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12857[13:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11957[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ac)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12882[13:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12522[13:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11537[13:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12727[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d) || (r_sys_run_step==9'h49)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10967[13:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11937[13:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12577[13:0] );

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12317[13:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12477[13:0] );

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12417[13:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12502[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10756[13:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11447[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12842[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12852[13:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11412[13:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11977[13:0] );

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12507[13:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12197[13:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11472[13:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11767[13:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11597[13:0] );

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12422[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11202[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10750[13:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12127[13:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12397[13:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12327[13:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12017[13:0] );

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11747[13:0] );

									end
									else
									if((r_sys_run_step==9'h30) || (r_sys_run_step==9'h4c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10982[13:0] );

									end
									else
									if((r_sys_run_step==9'h157)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12457[13:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11297[13:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11382[13:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11292[13:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12192[13:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12622[13:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11557[13:0] );

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11922[13:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11387[13:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12107[13:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12437[13:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12467[13:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11857[13:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11722[13:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11172[13:0] );

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12572[13:0] );

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12262[13:0] );

									end
									else
									if((r_sys_run_step==9'h183)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12677[13:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12227[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10762[13:0] );

									end
									else
									if((r_sys_run_step==9'h19c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12802[13:0] );

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11607[13:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11907[13:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11657[13:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12082[13:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12582[13:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12217[13:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12282[13:0] );

									end
									else
									if((r_sys_run_step==9'h199)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12787[13:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12222[13:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12352[13:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12377[13:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11792[13:0] );

									end
									else
									if((r_sys_run_step==9'h184)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12682[13:0] );

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12712[13:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12387[13:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11527[13:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11852[13:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12002[13:0] );

									end
									else
									if((r_sys_run_step==9'h12d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12247[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12922[13:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11987[13:0] );

									end
									else
									if((r_sys_run_step==9'h1af)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12897[13:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12172[13:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11467[13:0] );

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12602[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11247[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12847[13:0] );

									end
									else
									if((r_sys_run_step==9'h192)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12752[13:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11442[13:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12012[13:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11182[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12932[13:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12077[13:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11342[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a) || (r_sys_run_step==9'h46)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10952[13:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11402[13:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11457[13:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12512[13:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11692[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11167[13:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12187[13:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12742[13:0] );

									end
									else
									if((r_sys_run_step==9'hb) || (r_sys_run_step==9'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10786[13:0] );

									end
									else
									if((r_sys_run_step==9'h19e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12812[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11227[13:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11802[13:0] );

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12707[13:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12642[13:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11397[13:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12692[13:0] );

									end
									else
									if((r_sys_run_step==9'h35) || (r_sys_run_step==9'h51)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11007[13:0] );

									end
									else
									if((r_sys_run_step==9'h25) || (r_sys_run_step==9'h41)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10927[13:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11967[13:0] );

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12242[13:0] );

									end
									else
									if((r_sys_run_step==9'h31) || (r_sys_run_step==9'h4d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10987[13:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12732[13:0] );

									end
									else
									if((r_sys_run_step==9'h9) || (r_sys_run_step==9'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10774[13:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11352[13:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11322[13:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11627[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11222[13:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11982[13:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11392[13:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12232[13:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12392[13:0] );

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11752[13:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12067[13:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11542[13:0] );

									end
									else
									if((r_sys_run_step==9'h181)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12667[13:0] );

									end
									else
									if((r_sys_run_step==9'h10) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h3a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10816[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11187[13:0] );

									end
									else
									if((r_sys_run_step==9'h19a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12792[13:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12072[13:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11482[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11237[13:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12737[13:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11872[13:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11807[13:0] );

									end
									else
									if((r_sys_run_step==9'h12e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12252[13:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12662[13:0] );

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12762[13:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12632[13:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11577[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b) || (r_sys_run_step==9'h47)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10957[13:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11517[13:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11897[13:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12552[13:0] );

									end
									else
									if((r_sys_run_step==9'h2c) || (r_sys_run_step==9'h48)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10962[13:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12547[13:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12342[13:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12052[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12867[13:0] );

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12432[13:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12287[13:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11677[13:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12102[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10744[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11212[13:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12687[13:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11662[13:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11742[13:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11727[13:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12357[13:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12657[13:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11337[13:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12722[13:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12047[13:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11667[13:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11612[13:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12177[13:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12167[13:0] );

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12697[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11242[13:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12367[13:0] );

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11912[13:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12272[13:0] );

									end
									else
									if((r_sys_run_step==9'h11) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10822[13:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12302[13:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11952[13:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12092[13:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11637[13:0] );

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12137[13:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12007[13:0] );

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12257[13:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11647[13:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11307[13:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11882[13:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11487[13:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11587[13:0] );

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12142[13:0] );

									end
									else
									if((r_sys_run_step==9'heb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11917[13:0] );

									end
									else
									if((r_sys_run_step==9'hf) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10810[13:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12212[13:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12332[13:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11832[13:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12087[13:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11562[13:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12297[13:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12402[13:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11507[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11277[13:0] );

									end
									else
									if((r_sys_run_step==9'h67) || (r_sys_run_step==9'h68)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11257[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12917[13:0] );

									end
									else
									if((r_sys_run_step==9'h34) || (r_sys_run_step==9'h50)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11002[13:0] );

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11712[13:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11632[13:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12292[13:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12757[13:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12517[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e) || (r_sys_run_step==9'h4a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10972[13:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11972[13:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11932[13:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11672[13:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12637[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11252[13:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11452[13:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11797[13:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12347[13:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12497[13:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12487[13:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12132[13:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11942[13:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11312[13:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11787[13:0] );

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11497[13:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12472[13:0] );

									end
									else
									if((r_sys_run_step==9'h24) || (r_sys_run_step==9'h40)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10922[13:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12312[13:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12407[13:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12117[13:0] );

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12597[13:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12482[13:0] );

									end
									else
									if((r_sys_run_step==9'ha) || (r_sys_run_step==9'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10780[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12902[13:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11822[13:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12412[13:0] );

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12037[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11217[13:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11532[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ad)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12887[13:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12542[13:0] );

									end
									else
									if((r_sys_run_step==9'he) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10804[13:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12492[13:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12717[13:0] );

									end
									else
									if((r_sys_run_step==9'h36) || (r_sys_run_step==9'h52)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11012[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12827[13:0] );

									end
									else
									if((r_sys_run_step==9'h37) || (r_sys_run_step==9'h53)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11017[13:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11437[13:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11947[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11197[13:0] );

									end
									else
									if((r_sys_run_step==9'h171)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12587[13:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11732[13:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12372[13:0] );

									end
									else
									if((r_sys_run_step==9'h172)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12592[13:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12647[13:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11682[13:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11827[13:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11492[13:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12322[13:0] );

									end
									else
									if((r_sys_run_step==9'h8) || (r_sys_run_step==9'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10768[13:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11862[13:0] );

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12057[13:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12182[13:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11902[13:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11837[13:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11782[13:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11407[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11162[13:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12122[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ab)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12877[13:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11707[13:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12097[13:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11602[13:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11772[13:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12112[13:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11567[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12947[13:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11357[13:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12337[13:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11847[13:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12362[13:0] );

									end
									else
									if((r_sys_run_step==9'h182)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12672[13:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11817[13:0] );

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12032[13:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11687[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f) || (r_sys_run_step==9'h4b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10977[13:0] );

									end
									else
									if((r_sys_run_step==9'h33) || (r_sys_run_step==9'h4f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp10997[13:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12607[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11192[13:0] );

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12237[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12832[13:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12267[13:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11332[13:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12202[13:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11427[13:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11462[13:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11812[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12907[13:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12612[13:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11717[13:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11552[13:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11892[13:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11347[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12912[13:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12627[13:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12527[13:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12042[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12837[13:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12207[13:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11372[13:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11962[13:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12532[13:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11842[13:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11642[13:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11377[13:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11737[13:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12062[13:0] );

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12452[13:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12147[13:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11617[13:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11592[13:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11697[13:0] );

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12557[13:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp11997[13:0] );

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13308[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13263[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13438[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13268[13:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13403[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13423[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13208[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13318[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13133[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13243[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13138[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13193[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13228[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13313[13:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13298[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13048[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13303[13:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13083[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13108[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13358[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13128[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13333[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13203[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13463[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13000[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13418[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13273[13:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13293[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12988[13:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13408[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13113[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13258[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13088[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13173[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13383[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13353[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13148[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13363[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13238[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13338[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12982[13:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13188[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13158[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12994[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13343[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13393[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13036[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13078[13:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13072[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13198[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12964[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13373[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13118[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13042[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13006[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13278[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13323[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13153[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13218[13:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13398[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13060[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13030[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13018[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13123[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13283[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13054[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13328[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13163[13:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13288[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13143[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12976[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13443[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13448[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13024[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13428[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13098[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13453[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13178[13:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13066[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13458[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13348[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13253[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13103[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13368[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13378[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12970[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13223[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13168[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13012[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13183[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13468[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13233[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13413[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13433[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13213[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13388[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13093[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp12958[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp13248[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp7064;

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp7069;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h27)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp7082;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp7329;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp295_float;

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp242_float;

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp304_float;

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp193_float;

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp177_float;

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp246_float;

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp198_float;

									end
									else
									if((r_sys_run_step==9'h27) || (r_sys_run_step==9'h5d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp380_float;

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp95_float;

									end
									else
									if((r_sys_run_step==9'h1a) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h64)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp387_float;

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp133_float;

									end
									else
									if((r_sys_run_step==9'h1b9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp136_float;

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp144_float;

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp319_float;

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp128_float;

									end
									else
									if((r_sys_run_step==9'h19c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp201_float;

									end
									else
									if((r_sys_run_step==9'h184)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp274_float;

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp186_float;

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp117_float;

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp155_float;

									end
									else
									if((r_sys_run_step==9'h1aa)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp300_float;

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp370_float;

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp110_float;

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp161_float;

									end
									else
									if((r_sys_run_step==9'h19d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp175_float;

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp159_float;

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp91_float;

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp351_float;

									end
									else
									if((r_sys_run_step==9'h183)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp289_float;

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp249_float;

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp78_float;

									end
									else
									if((r_sys_run_step==9'h1a4)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==9'h22) || (r_sys_run_step==9'h36)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp373_float;

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp199_float;

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp122_float;

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp306_float;

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp82_float;

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp344_float;

									end
									else
									if((r_sys_run_step==9'h1b1)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp176_float;

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp124_float;

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp81_float;

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp297_float;

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp205_float;

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp220_float;

									end
									else
									if((r_sys_run_step==9'h196)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp312_float;

									end
									else
									if((r_sys_run_step==9'h17) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h61)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp390_float;

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp247_float;

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp286_float;

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp243_float;

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp361_float;

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp283_float;

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp342_float;

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp268_float;

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp231_float;

									end
									else
									if((r_sys_run_step==9'h1ad)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp251_float;

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp332_float;

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp261_float;

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp318_float;

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp280_float;

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp194_float;

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp347_float;

									end
									else
									if((r_sys_run_step==9'h1d) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h67)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp384_float;

									end
									else
									if((r_sys_run_step==9'h1ae)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp239_float;

									end
									else
									if((r_sys_run_step==9'h19a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp238_float;

									end
									else
									if((r_sys_run_step==9'h26) || (r_sys_run_step==9'h5c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp381_float;

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp343_float;

									end
									else
									if((r_sys_run_step==9'h171)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp252_float;

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp211_float;

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp271_float;

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp216_float;

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp142_float;

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp140_float;

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp301_float;

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp290_float;

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp180_float;

									end
									else
									if((r_sys_run_step==9'h25) || (r_sys_run_step==9'h5b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp382_float;

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp123_float;

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp62_float;

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp320_float;

									end
									else
									if((r_sys_run_step==9'h1b3)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp152_float;

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==9'h23) || (r_sys_run_step==9'h37)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp372_float;

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp294_float;

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp352_float;

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp241_float;

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp340_float;

									end
									else
									if((r_sys_run_step==9'h1ab)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp288_float;

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp282_float;

									end
									else
									if((r_sys_run_step==9'h16) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h60)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp391_float;

									end
									else
									if((r_sys_run_step==9'h1a3)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp132_float;

									end
									else
									if((r_sys_run_step==9'h1b) || (r_sys_run_step==9'h2f) || (r_sys_run_step==9'h65)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp386_float;

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp116_float;

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp292_float;

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp187_float;

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp77_float;

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==9'h157)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp358_float;

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp98_float;

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp74_float;

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp356_float;

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp284_float;

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp260_float;

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp141_float;

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp94_float;

									end
									else
									if((r_sys_run_step==9'h1a7)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp360_float;

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp210_float;

									end
									else
									if((r_sys_run_step==9'h1b2)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp165_float;

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp367_float;

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==9'h19) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h63)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp388_float;

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp223_float;

									end
									else
									if((r_sys_run_step==9'h1b4)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp126_float;

									end
									else
									if((r_sys_run_step==9'h195)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp323_float;

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp139_float;

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp354_float;

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp310_float;

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp230_float;

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp258_float;

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp307_float;

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp226_float;

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp169_float;

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp285_float;

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp219_float;

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp119_float;

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp120_float;

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp192_float;

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp259_float;

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp311_float;

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp108_float;

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp267_float;

									end
									else
									if((r_sys_run_step==9'h1a8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp348_float;

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp88_float;

									end
									else
									if((r_sys_run_step==9'h29) || (r_sys_run_step==9'h5f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp378_float;

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp168_float;

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==9'h1a2)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp99_float;

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp87_float;

									end
									else
									if((r_sys_run_step==9'h199)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp250_float;

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp173_float;

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp147_float;

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp190_float;

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp235_float;

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp206_float;

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==9'h19e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp163_float;

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp83_float;

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp305_float;

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp273_float;

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp80_float;

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp293_float;

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp363_float;

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp121_float;

									end
									else
									if((r_sys_run_step==9'h12d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp309_float;

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp195_float;

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp303_float;

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp266_float;

									end
									else
									if((r_sys_run_step==9'h188)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp200_float;

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp151_float;

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp255_float;

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp204_float;

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp334_float;

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp264_float;

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp257_float;

									end
									else
									if((r_sys_run_step==9'h19b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp225_float;

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp355_float;

									end
									else
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h15)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp10734;

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp365_float;

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp149_float;

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp115_float;

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp138_float;

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp222_float;

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp331_float;

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp281_float;

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp197_float;

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp253_float;

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp90_float;

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp135_float;

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp302_float;

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp191_float;

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp234_float;

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp146_float;

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp364_float;

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp162_float;

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp102_float;

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp330_float;

									end
									else
									if((r_sys_run_step==9'h1a0)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp125_float;

									end
									else
									if((r_sys_run_step==9'h19f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp150_float;

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp321_float;

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp97_float;

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp335_float;

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp338_float;

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp214_float;

									end
									else
									if((r_sys_run_step==9'h1b5)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp113_float;

									end
									else
									if((r_sys_run_step==9'h192)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==9'h24) || (r_sys_run_step==9'h5a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp383_float;

									end
									else
									if((r_sys_run_step==9'h1b8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp137_float;

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp229_float;

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp111_float;

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp296_float;

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp328_float;

									end
									else
									if((r_sys_run_step==9'h1b7)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp75_float;

									end
									else
									if((r_sys_run_step==9'h1b6)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp101_float;

									end
									else
									if((r_sys_run_step==9'heb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp188_float;

									end
									else
									if((r_sys_run_step==9'h1a1)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp112_float;

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp217_float;

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp76_float;

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp209_float;

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp208_float;

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp184_float;

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp118_float;

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp100_float;

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp160_float;

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp244_float;

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp215_float;

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp237_float;

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp167_float;

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp346_float;

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp333_float;

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp329_float;

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp179_float;

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp298_float;

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp369_float;

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp314_float;

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp183_float;

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp181_float;

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp322_float;

									end
									else
									if((r_sys_run_step==9'h12e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==9'h181)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp325_float;

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp164_float;

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp106_float;

									end
									else
									if((r_sys_run_step==9'h198)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp275_float;

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp131_float;

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp359_float;

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp345_float;

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp104_float;

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp158_float;

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp218_float;

									end
									else
									if((r_sys_run_step==9'h172)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp236_float;

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp114_float;

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp130_float;

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp353_float;

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp156_float;

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp339_float;

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==9'h197)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp287_float;

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp263_float;

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp291_float;

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp154_float;

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp262_float;

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp265_float;

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp277_float;

									end
									else
									if((r_sys_run_step==9'h1a6)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp316_float;

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp349_float;

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp336_float;

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp254_float;

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp233_float;

									end
									else
									if((r_sys_run_step==9'h28) || (r_sys_run_step==9'h5e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp379_float;

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp270_float;

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp245_float;

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp109_float;

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp92_float;

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp93_float;

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp341_float;

									end
									else
									if((r_sys_run_step==9'h1a5)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp178_float;

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp157_float;

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp337_float;

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp170_float;

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp357_float;

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp143_float;

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp279_float;

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp228_float;

									end
									else
									if((r_sys_run_step==9'h1f) || (r_sys_run_step==9'h33)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp376_float;

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp317_float;

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp366_float;

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp96_float;

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp256_float;

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp350_float;

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp84_float;

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp371_float;

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp196_float;

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp248_float;

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp185_float;

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp315_float;

									end
									else
									if((r_sys_run_step==9'h20) || (r_sys_run_step==9'h34)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp375_float;

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp134_float;

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==9'h18) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h62)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp389_float;

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp299_float;

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp145_float;

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp172_float;

									end
									else
									if((r_sys_run_step==9'h21) || (r_sys_run_step==9'h35)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp374_float;

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp278_float;

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp148_float;

									end
									else
									if((r_sys_run_step==9'h1ac)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp276_float;

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp129_float;

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp89_float;

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp103_float;

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp207_float;

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp166_float;

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp189_float;

									end
									else
									if((r_sys_run_step==9'h1b0)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp202_float;

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==9'h1af)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp227_float;

									end
									else
									if((r_sys_run_step==9'h1c) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h66)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp385_float;

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp221_float;

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp174_float;

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp272_float;

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp171_float;

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp212_float;

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp127_float;

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp153_float;

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp213_float;

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp232_float;

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp182_float;

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp368_float;

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp308_float;

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp326_float;

									end
									else
									if((r_sys_run_step==9'h1a9)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp324_float;

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp203_float;

									end
									else
									if((r_sys_run_step==9'h182)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp313_float;

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp240_float;

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp269_float;

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp85_float;

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp105_float;

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp362_float;

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==9'h1e) || (r_sys_run_step==9'h32)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp377_float;

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp224_float;

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp327_float;

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp107_float;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h56)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp75_float;

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp58_float;

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp82_float;

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp81_float;

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp72_float;

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp60_float;

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp89_float;

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp76_float;

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp70_float;

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp51_float;

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp95_float;

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp59_float;

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp73_float;

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp65_float;

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp92_float;

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp93_float;

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp77_float;

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp53_float;

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp74_float;

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp54_float;

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp66_float;

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp90_float;

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp71_float;

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp88_float;

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp64_float;

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp86_float;

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp87_float;

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp67_float;

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp52_float;

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp79_float;

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp48_float;

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp94_float;

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp68_float;

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp102_float;

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp84_float;

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp91_float;

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp63_float;

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp78_float;

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp61_float;

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp83_float;

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp85_float;

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp57_float;

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp49_float;

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp80_float;

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp62_float;

									end
									else
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h15)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp12960;

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp50_float;

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp69_float;

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp56_float;

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp55_float;

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp23_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h3)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h27)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1b3)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6c)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h1b9)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h64)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp27[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h3d) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h41) || (9'h43<=r_sys_run_step && r_sys_run_step<=9'h47)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp32[13:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1889[13:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3089[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1793[13:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2105[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp881[13:0] );

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4649[13:0] );

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3977[13:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3869[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp677[13:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4565[13:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1961[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1781[13:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1997[13:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3221[13:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4757[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp665[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp785[13:0] );

									end
									else
									if((r_sys_run_step==9'h15) || (r_sys_run_step==9'h17)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp845[13:0] );

									end
									else
									if((r_sys_run_step==9'h192)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5417[13:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4793[13:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4265[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1805[13:0] );

									end
									else
									if((r_sys_run_step==9'heb) || (r_sys_run_step==9'hec)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3413[13:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3509[13:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2597[13:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4721[13:0] );

									end
									else
									if((r_sys_run_step==9'h19f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5573[13:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5357[13:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5201[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ac)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5729[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1661[13:0] );

									end
									else
									if((r_sys_run_step==9'h19b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5525[13:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2117[13:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3209[13:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4133[13:0] );

									end
									else
									if((r_sys_run_step==9'h1aa)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5705[13:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2993[13:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3449[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp773[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp713[13:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4157[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1289[13:0] );

									end
									else
									if((r_sys_run_step==9'h80) || (r_sys_run_step==9'h81)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2129[13:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2369[13:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3245[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1253[13:0] );

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5321[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1241[13:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2873[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1493[13:0] );

									end
									else
									if((r_sys_run_step==9'hc1) || (r_sys_run_step==9'hc3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2909[13:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2681[13:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2633[13:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4685[13:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3305[13:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4097[13:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4841[13:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3533[13:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2801[13:0] );

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3437[13:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4673[13:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2945[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1577[13:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3725[13:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5009[13:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2789[13:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4577[13:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2249[13:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3833[13:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3473[13:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4817[13:0] );

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5045[13:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2765[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1841[13:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2717[13:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1973[13:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5345[13:0] );

									end
									else
									if((r_sys_run_step==9'h96) || (r_sys_run_step==9'h98)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2393[13:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5381[13:0] );

									end
									else
									if((r_sys_run_step==9'h197) || (r_sys_run_step==9'h199)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5477[13:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5117[13:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2693[13:0] );

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5309[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ad)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5741[13:0] );

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5057[13:0] );

									end
									else
									if((r_sys_run_step==9'h172)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5033[13:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2021[13:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4337[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp929[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1769[13:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2861[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1397[13:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4013[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1853[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1457[13:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4457[13:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4505[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1733[13:0] );

									end
									else
									if((r_sys_run_step==9'h117) || (r_sys_run_step==9'h118)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3941[13:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2489[13:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4445[13:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2513[13:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2321[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp629[13:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3557[13:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3629[13:0] );

									end
									else
									if((r_sys_run_step==9'h19d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5549[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1001[13:0] );

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3017[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp989[13:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2825[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1757[13:0] );

									end
									else
									if((r_sys_run_step==9'h12b) || (r_sys_run_step==9'h12d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4181[13:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2453[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1589[13:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2837[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1217[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp941[13:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2981[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1469[13:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2045[13:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3461[13:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1937[13:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1925[13:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2213[13:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3617[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1565[13:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4925[13:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1385[13:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4169[13:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3881[13:0] );

									end
									else
									if((r_sys_run_step==9'h156) || (r_sys_run_step==9'h157)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4697[13:0] );

									end
									else
									if((r_sys_run_step==9'h19e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5561[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp905[13:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3713[13:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3845[13:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3929[13:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5273[13:0] );

									end
									else
									if((r_sys_run_step==9'h196)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5465[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1313[13:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3857[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5693[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1073[13:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4145[13:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4853[13:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2777[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp893[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1481[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1181[13:0] );

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5405[13:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3269[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp917[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp641[13:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3329[13:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3641[13:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4913[13:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5429[13:0] );

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4001[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1865[13:0] );

									end
									else
									if((r_sys_run_step==9'h19c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5537[13:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3257[13:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2885[13:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3233[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1829[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1109[13:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2273[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1445[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1709[13:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3809[13:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4025[13:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2525[13:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4865[13:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3389[13:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2753[13:0] );

									end
									else
									if((r_sys_run_step==9'hc0) || (r_sys_run_step==9'hc2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2897[13:0] );

									end
									else
									if((r_sys_run_step==9'h188)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5297[13:0] );

									end
									else
									if((r_sys_run_step==9'h16b) || (r_sys_run_step==9'h16d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4949[13:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2645[13:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4889[13:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4325[13:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2849[13:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4541[13:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2081[13:0] );

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4241[13:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2429[13:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2285[13:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3653[13:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3065[13:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3353[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5669[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5633[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1673[13:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4049[13:0] );

									end
									else
									if((r_sys_run_step==9'h101) || (r_sys_run_step==9'h103)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3677[13:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2225[13:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2465[13:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1985[13:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3137[13:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2165[13:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4481[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1409[13:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2621[13:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3125[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1433[13:0] );

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3005[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp749[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5621[13:0] );

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3401[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1169[13:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2057[13:0] );

									end
									else
									if((r_sys_run_step==9'h95) || (r_sys_run_step==9'h97)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2381[13:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5189[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1097[13:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4517[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp725[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp605[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp761[13:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3317[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1745[13:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4277[13:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2705[13:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4769[13:0] );

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4229[13:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3101[13:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1913[13:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5261[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1049[13:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4073[13:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2561[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp797[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp965[13:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2189[13:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2033[13:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3293[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1277[13:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1949[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp617[13:0] );

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4613[13:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5093[13:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5393[13:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4589[13:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3341[13:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3281[13:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3965[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5597[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1085[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1157[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1421[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5645[13:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3197[13:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2441[13:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4409[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1901[13:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3581[13:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3185[13:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4289[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1553[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1145[13:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4397[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp821[13:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4997[13:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3905[13:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4061[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1349[13:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4901[13:0] );

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4625[13:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5141[13:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2813[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1193[13:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3773[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1697[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1265[13:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2153[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1337[13:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3521[13:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4601[13:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3077[13:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3161[13:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3053[13:0] );

									end
									else
									if((r_sys_run_step==9'h198) || (r_sys_run_step==9'h19a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5489[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1205[13:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3485[13:0] );

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4637[13:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3377[13:0] );

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3029[13:0] );

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4829[13:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3497[13:0] );

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5441[13:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4301[13:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4361[13:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3785[13:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4037[13:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5153[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp653[13:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2093[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1505[13:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3173[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp689[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1025[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5609[13:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4385[13:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2009[13:0] );

									end
									else
									if((r_sys_run_step==9'h195)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5453[13:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2969[13:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4745[13:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2357[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1517[13:0] );

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5285[13:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4109[13:0] );

									end
									else
									if((r_sys_run_step==9'h55) || (r_sys_run_step==9'h57)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1613[13:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2729[13:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2261[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1529[13:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5069[13:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3737[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp977[13:0] );

									end
									else
									if((r_sys_run_step==9'h16c) || (r_sys_run_step==9'h16e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4961[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1037[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp701[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1325[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1061[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp953[13:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2573[13:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4433[13:0] );

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3749[13:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2501[13:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3989[13:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2741[13:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5165[13:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4781[13:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2537[13:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3605[13:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3917[13:0] );

									end
									else
									if((r_sys_run_step==9'h182) || (r_sys_run_step==9'h184)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5225[13:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2177[13:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4529[13:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3365[13:0] );

									end
									else
									if((r_sys_run_step==9'h100) || (r_sys_run_step==9'h102)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3665[13:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5129[13:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2201[13:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2237[13:0] );

									end
									else
									if((r_sys_run_step==9'h12c) || (r_sys_run_step==9'h12e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4193[13:0] );

									end
									else
									if((r_sys_run_step==9'h56) || (r_sys_run_step==9'h58)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1625[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1817[13:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4085[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1301[13:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4313[13:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5105[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1229[13:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5081[13:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4553[13:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3821[13:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2957[13:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3113[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5657[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ab)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5717[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5681[13:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4733[13:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3149[13:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4661[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp737[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1721[13:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2549[13:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4805[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1541[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1877[13:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4877[13:0] );

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4373[13:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2333[13:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5369[13:0] );

									end
									else
									if((r_sys_run_step==9'h171)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5021[13:0] );

									end
									else
									if((r_sys_run_step==9'h14) || (r_sys_run_step==9'h16)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp833[13:0] );

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2585[13:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3569[13:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2477[13:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2309[13:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3545[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5585[13:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3893[13:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4469[13:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2297[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp593[13:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4349[13:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3041[13:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5333[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1685[13:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2609[13:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4421[13:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3761[13:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4937[13:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4253[13:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2345[13:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3797[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1013[13:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2069[13:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4493[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp809[13:0] );

									end
									else
									if((r_sys_run_step==9'h40) || (r_sys_run_step==9'h41)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1361[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1601[13:0] );

									end
									else
									if((r_sys_run_step==9'hac) || (r_sys_run_step==9'had)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp2657[13:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5177[13:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp4121[13:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp3593[13:0] );

									end
									else
									if((r_sys_run_step==9'h181) || (r_sys_run_step==9'h183)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5213[13:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h25)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6203[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6383[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6311[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6491[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6911[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5867[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6395[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6875[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5795[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6719[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5963[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6959[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6923[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6635[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5903[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6059[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6899[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6671[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6215[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6179[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6647[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6839[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5879[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6947[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5987[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6119[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6431[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6575[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5783[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6683[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6167[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6263[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5759[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6863[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6971[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6371[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6755[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6047[13:0] );

									end
									else
									if((r_sys_run_step==9'h56) || (r_sys_run_step==9'h58)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6791[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5951[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6983[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6611[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6503[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6023[13:0] );

									end
									else
									if((r_sys_run_step==9'h55) || (r_sys_run_step==9'h57)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6779[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6131[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6731[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp7019[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6419[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp7007[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f) || (r_sys_run_step==9'h41)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6515[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5855[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6455[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6083[13:0] );

									end
									else
									if((r_sys_run_step==9'h14) || (r_sys_run_step==9'h15)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5999[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6743[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6767[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6155[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6599[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6887[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6239[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5831[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6443[13:0] );

									end
									else
									if((r_sys_run_step==9'h29) || (r_sys_run_step==9'h2b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6251[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6299[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5915[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6467[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5819[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6479[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6107[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6659[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6095[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5891[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp7043[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6587[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6347[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6335[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5807[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6191[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6563[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp7031[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6707[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6143[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6227[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6323[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6995[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5771[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5843[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5939[13:0] );

									end
									else
									if((r_sys_run_step==9'h40) || (r_sys_run_step==9'h42)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6527[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6827[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6359[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6695[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6407[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6935[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6071[13:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6035[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5975[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6623[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp5927[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp6851[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h3d) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h41) || (9'h43<=r_sys_run_step && r_sys_run_step<=9'h47)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h3d) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h41) || (9'h43<=r_sys_run_step && r_sys_run_step<=9'h47)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1ad)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6b)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_addr_1 <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp41[13:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1889[13:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3089[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1793[13:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2105[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp881[13:0] );

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4649[13:0] );

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3977[13:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3869[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp677[13:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4565[13:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1961[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1781[13:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1997[13:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3221[13:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4757[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp665[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp785[13:0] );

									end
									else
									if((r_sys_run_step==9'h15) || (r_sys_run_step==9'h17)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp845[13:0] );

									end
									else
									if((r_sys_run_step==9'h192)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5417[13:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4793[13:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4265[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1805[13:0] );

									end
									else
									if((r_sys_run_step==9'heb) || (r_sys_run_step==9'hec)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3413[13:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3509[13:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2597[13:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4721[13:0] );

									end
									else
									if((r_sys_run_step==9'h19f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5573[13:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5357[13:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5201[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ac)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5729[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1661[13:0] );

									end
									else
									if((r_sys_run_step==9'h19b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5525[13:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2117[13:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3209[13:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4133[13:0] );

									end
									else
									if((r_sys_run_step==9'h1aa)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5705[13:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2993[13:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3449[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp773[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp713[13:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4157[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1289[13:0] );

									end
									else
									if((r_sys_run_step==9'h80) || (r_sys_run_step==9'h81)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2129[13:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2369[13:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3245[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1253[13:0] );

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5321[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1241[13:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2873[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1493[13:0] );

									end
									else
									if((r_sys_run_step==9'hc1) || (r_sys_run_step==9'hc3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2909[13:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2681[13:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2633[13:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4685[13:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3305[13:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4097[13:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4841[13:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3533[13:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2801[13:0] );

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3437[13:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4673[13:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2945[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1577[13:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3725[13:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5009[13:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2789[13:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4577[13:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2249[13:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3833[13:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3473[13:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4817[13:0] );

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5045[13:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2765[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1841[13:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2717[13:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1973[13:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5345[13:0] );

									end
									else
									if((r_sys_run_step==9'h96) || (r_sys_run_step==9'h98)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2393[13:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5381[13:0] );

									end
									else
									if((r_sys_run_step==9'h197) || (r_sys_run_step==9'h199)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5477[13:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5117[13:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2693[13:0] );

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5309[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ad)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5741[13:0] );

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5057[13:0] );

									end
									else
									if((r_sys_run_step==9'h172)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5033[13:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2021[13:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4337[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp929[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1769[13:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2861[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1397[13:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4013[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1853[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1457[13:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4457[13:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4505[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1733[13:0] );

									end
									else
									if((r_sys_run_step==9'h117) || (r_sys_run_step==9'h118)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3941[13:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2489[13:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4445[13:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2513[13:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2321[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp629[13:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3557[13:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3629[13:0] );

									end
									else
									if((r_sys_run_step==9'h19d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5549[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1001[13:0] );

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3017[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp989[13:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2825[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1757[13:0] );

									end
									else
									if((r_sys_run_step==9'h12b) || (r_sys_run_step==9'h12d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4181[13:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2453[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1589[13:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2837[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1217[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp941[13:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2981[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1469[13:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2045[13:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3461[13:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1937[13:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1925[13:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2213[13:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3617[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1565[13:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4925[13:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1385[13:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4169[13:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3881[13:0] );

									end
									else
									if((r_sys_run_step==9'h156) || (r_sys_run_step==9'h157)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4697[13:0] );

									end
									else
									if((r_sys_run_step==9'h19e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5561[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp905[13:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3713[13:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3845[13:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3929[13:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5273[13:0] );

									end
									else
									if((r_sys_run_step==9'h196)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5465[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1313[13:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3857[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5693[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1073[13:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4145[13:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4853[13:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2777[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp893[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1481[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1181[13:0] );

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5405[13:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3269[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp917[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp641[13:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3329[13:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3641[13:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4913[13:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5429[13:0] );

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4001[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1865[13:0] );

									end
									else
									if((r_sys_run_step==9'h19c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5537[13:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3257[13:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2885[13:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3233[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1829[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1109[13:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2273[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1445[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1709[13:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3809[13:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4025[13:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2525[13:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4865[13:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3389[13:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2753[13:0] );

									end
									else
									if((r_sys_run_step==9'hc0) || (r_sys_run_step==9'hc2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2897[13:0] );

									end
									else
									if((r_sys_run_step==9'h188)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5297[13:0] );

									end
									else
									if((r_sys_run_step==9'h16b) || (r_sys_run_step==9'h16d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4949[13:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2645[13:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4889[13:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4325[13:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2849[13:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4541[13:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2081[13:0] );

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4241[13:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2429[13:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2285[13:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3653[13:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3065[13:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3353[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5669[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5633[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1673[13:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4049[13:0] );

									end
									else
									if((r_sys_run_step==9'h101) || (r_sys_run_step==9'h103)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3677[13:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2225[13:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2465[13:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1985[13:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3137[13:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2165[13:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4481[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1409[13:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2621[13:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3125[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1433[13:0] );

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3005[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp749[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5621[13:0] );

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3401[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1169[13:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2057[13:0] );

									end
									else
									if((r_sys_run_step==9'h95) || (r_sys_run_step==9'h97)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2381[13:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5189[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1097[13:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4517[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp725[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp605[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp761[13:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3317[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1745[13:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4277[13:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2705[13:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4769[13:0] );

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4229[13:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3101[13:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1913[13:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5261[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1049[13:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4073[13:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2561[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp797[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp965[13:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2189[13:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2033[13:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3293[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1277[13:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1949[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp617[13:0] );

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4613[13:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5093[13:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5393[13:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4589[13:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3341[13:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3281[13:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3965[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5597[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1085[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1157[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1421[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5645[13:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3197[13:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2441[13:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4409[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1901[13:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3581[13:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3185[13:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4289[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1553[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1145[13:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4397[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp821[13:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4997[13:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3905[13:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4061[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1349[13:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4901[13:0] );

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4625[13:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5141[13:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2813[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1193[13:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3773[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1697[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1265[13:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2153[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1337[13:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3521[13:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4601[13:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3077[13:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3161[13:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3053[13:0] );

									end
									else
									if((r_sys_run_step==9'h198) || (r_sys_run_step==9'h19a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5489[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1205[13:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3485[13:0] );

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4637[13:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3377[13:0] );

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3029[13:0] );

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4829[13:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3497[13:0] );

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5441[13:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4301[13:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4361[13:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3785[13:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4037[13:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5153[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp653[13:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2093[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1505[13:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3173[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp689[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1025[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5609[13:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4385[13:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2009[13:0] );

									end
									else
									if((r_sys_run_step==9'h195)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5453[13:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2969[13:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4745[13:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2357[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1517[13:0] );

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5285[13:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4109[13:0] );

									end
									else
									if((r_sys_run_step==9'h55) || (r_sys_run_step==9'h57)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1613[13:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2729[13:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2261[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1529[13:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5069[13:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3737[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp977[13:0] );

									end
									else
									if((r_sys_run_step==9'h16c) || (r_sys_run_step==9'h16e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4961[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1037[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp701[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1325[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1061[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp953[13:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2573[13:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4433[13:0] );

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3749[13:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2501[13:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3989[13:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2741[13:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5165[13:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4781[13:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2537[13:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3605[13:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3917[13:0] );

									end
									else
									if((r_sys_run_step==9'h182) || (r_sys_run_step==9'h184)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5225[13:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2177[13:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4529[13:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3365[13:0] );

									end
									else
									if((r_sys_run_step==9'h100) || (r_sys_run_step==9'h102)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3665[13:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5129[13:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2201[13:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2237[13:0] );

									end
									else
									if((r_sys_run_step==9'h12c) || (r_sys_run_step==9'h12e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4193[13:0] );

									end
									else
									if((r_sys_run_step==9'h56) || (r_sys_run_step==9'h58)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1625[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1817[13:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4085[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1301[13:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4313[13:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5105[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1229[13:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5081[13:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4553[13:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3821[13:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2957[13:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3113[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5657[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ab)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5717[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5681[13:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4733[13:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3149[13:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4661[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp737[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1721[13:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2549[13:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4805[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1541[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1877[13:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4877[13:0] );

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4373[13:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2333[13:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5369[13:0] );

									end
									else
									if((r_sys_run_step==9'h171)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5021[13:0] );

									end
									else
									if((r_sys_run_step==9'h14) || (r_sys_run_step==9'h16)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp833[13:0] );

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2585[13:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3569[13:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2477[13:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2309[13:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3545[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5585[13:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3893[13:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4469[13:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2297[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp593[13:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4349[13:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3041[13:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5333[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1685[13:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2609[13:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4421[13:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3761[13:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4937[13:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4253[13:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2345[13:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3797[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1013[13:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2069[13:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4493[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp809[13:0] );

									end
									else
									if((r_sys_run_step==9'h40) || (r_sys_run_step==9'h41)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1361[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1601[13:0] );

									end
									else
									if((r_sys_run_step==9'hac) || (r_sys_run_step==9'had)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp2657[13:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5177[13:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp4121[13:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp3593[13:0] );

									end
									else
									if((r_sys_run_step==9'h181) || (r_sys_run_step==9'h183)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5213[13:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h25)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6203[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6383[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6311[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6491[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6911[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5867[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6395[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6875[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5795[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6719[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5963[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6959[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6923[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6635[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5903[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6059[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6899[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6671[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6215[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6179[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6647[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6839[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5879[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6947[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5987[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6119[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6431[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6575[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5783[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6683[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6167[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a) || (r_sys_run_step==9'h2c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6263[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5759[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6863[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6971[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6371[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6755[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6047[13:0] );

									end
									else
									if((r_sys_run_step==9'h56) || (r_sys_run_step==9'h58)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6791[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5951[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6983[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6611[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6503[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6023[13:0] );

									end
									else
									if((r_sys_run_step==9'h55) || (r_sys_run_step==9'h57)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6779[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6131[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6731[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp7019[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6419[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp7007[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f) || (r_sys_run_step==9'h41)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6515[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5855[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6455[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6083[13:0] );

									end
									else
									if((r_sys_run_step==9'h14) || (r_sys_run_step==9'h15)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5999[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6743[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6767[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6155[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6599[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6887[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6239[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5831[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6443[13:0] );

									end
									else
									if((r_sys_run_step==9'h29) || (r_sys_run_step==9'h2b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6251[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6299[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5915[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6467[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5819[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6479[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6107[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6659[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6095[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5891[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp7043[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6587[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6347[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6335[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5807[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6191[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6563[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp7031[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6707[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6143[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6227[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6323[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6995[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5771[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5843[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5939[13:0] );

									end
									else
									if((r_sys_run_step==9'h40) || (r_sys_run_step==9'h42)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6527[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6827[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6359[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6695[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6407[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6935[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6071[13:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6035[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5975[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6623[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp5927[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp6851[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_V_3_datain_1 <= w_sys_tmp25;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h1ad)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h6b)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_V_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_29 <= w_sys_tmp14;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1af)) begin
										r_run_k_29 <= w_sys_tmp5752;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_29 <= w_sys_tmp5753;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6d)) begin
										r_run_k_29 <= w_sys_tmp7054;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_run_k_29 <= w_sys_tmp7074;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_29 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b5)) begin
										r_run_k_29 <= w_sys_tmp10065;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_29 <= w_sys_tmp10066;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6e)) begin
										r_run_k_29 <= w_sys_tmp10725;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_29 <= w_sys_tmp10726;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b9)) begin
										r_run_k_29 <= w_sys_tmp12951;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_k_29 <= w_sys_tmp12952;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h64)) begin
										r_run_k_29 <= w_sys_tmp13472;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_30 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_run_j_30 <= w_sys_tmp48;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_j_30 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0) || (r_sys_run_step==9'h2) || (r_sys_run_step==9'h4) || (r_sys_run_step==9'h6) || (r_sys_run_step==9'h8) || (r_sys_run_step==9'ha) || (r_sys_run_step==9'hc) || (r_sys_run_step==9'he) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h14) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h26)) begin
										r_run_j_30 <= w_sys_tmp7089;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h25)) begin
										r_run_j_30 <= w_sys_tmp7318;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_run_j_30 <= w_sys_tmp7330;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_n_31 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_n_31 <= w_sys_tmp7057;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_mx_32 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_my_33 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_dt_34 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_dx_35 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_dy_36 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_r1_37 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_r2_38 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_r3_39 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_r4_40 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11) || (r_sys_run_step==9'h3b)) begin
										r_run_YY_41 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==9'h1e) || (r_sys_run_step==9'h27) || (r_sys_run_step==9'h30) || (r_sys_run_step==9'h37)) begin
										r_run_YY_41 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_run_YY_41 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_run_YY_41 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==9'h21) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h33) || (r_sys_run_step==9'h39)) begin
										r_run_YY_41 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==9'h15) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h35)) begin
										r_run_YY_41 <= r_sys_tmp14_float;

									end
									else
									if((r_sys_run_step==9'hc) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'he)) begin
										r_run_YY_41 <= w_sys_tmp18;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_kx_42 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_ky_43 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_nlast_44 <= w_sys_intOne;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_45 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_run_copy0_j_45 <= w_sys_tmp45;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy1_j_46 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h22) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h28) || (r_sys_run_step==9'h2b) || (r_sys_run_step==9'h2e) || (r_sys_run_step==9'h31) || (r_sys_run_step==9'h34) || (r_sys_run_step==9'h37) || (r_sys_run_step==9'h39) || (r_sys_run_step==9'h3b) || (r_sys_run_step==9'h3d) || (r_sys_run_step==9'h3f) || (r_sys_run_step==9'h41) || (9'h43<=r_sys_run_step && r_sys_run_step<=9'h47)) begin
										r_run_copy1_j_46 <= w_sys_tmp46;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy2_j_47 <= r_run_j_30;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_run_copy2_j_47 <= w_sys_tmp47;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_run_copy0_j_48 <= r_run_j_30;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1) || (r_sys_run_step==9'h3) || (r_sys_run_step==9'h5) || (r_sys_run_step==9'h7) || (r_sys_run_step==9'h9) || (r_sys_run_step==9'hb) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h17) || (r_sys_run_step==9'h19) || (r_sys_run_step==9'h1b) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h1f) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h25) || (r_sys_run_step==9'h27)) begin
										r_run_copy0_j_48 <= w_sys_tmp7088;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h13: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub19_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub19_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b4)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10054[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a1)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp9928[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a3)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp9952[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ab)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10000[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a7)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp9976[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a9)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp9988[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ad)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10012[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ae)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10018[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b1)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10036[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b5)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10060[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a4)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp9958[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a8)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp9982[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b3)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10048[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a6)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp9970[13:0] );

									end
									else
									if((r_sys_run_step==9'h1af)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10024[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a5)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp9964[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ac)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10006[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a2)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp9934[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b0)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10030[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b2)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp10042[13:0] );

									end
									else
									if((r_sys_run_step==9'h1aa)) begin
										r_sub19_T_addr <= $signed( w_sys_tmp9994[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h1a1<=r_sys_run_step && r_sys_run_step<=9'h1b5)) begin
										r_sub19_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h1a1<=r_sys_run_step && r_sys_run_step<=9'h1b5)) begin
										r_sub19_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a9)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5669[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a7)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5645[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a6)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5633[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a4)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5609[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ab)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5693[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a1)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5573[13:0] );

									end
									else
									if((r_sys_run_step==9'h19b)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5477[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a5)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5621[13:0] );

									end
									else
									if((r_sys_run_step==9'h19c)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5489[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ae)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5729[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a8)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5657[13:0] );

									end
									else
									if((r_sys_run_step==9'h19d)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5525[13:0] );

									end
									else
									if((r_sys_run_step==9'h19e)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5537[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ad)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5717[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a3)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5597[13:0] );

									end
									else
									if((r_sys_run_step==9'h1af)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5741[13:0] );

									end
									else
									if((r_sys_run_step==9'h1aa)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5681[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ac)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5705[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a0)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5561[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a2)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5585[13:0] );

									end
									else
									if((r_sys_run_step==9'h19f)) begin
										r_sub19_V_addr <= $signed( w_sys_tmp5549[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h19b<=r_sys_run_step && r_sys_run_step<=9'h1af)) begin
										r_sub19_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h19b<=r_sys_run_step && r_sys_run_step<=9'h1af)) begin
										r_sub19_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a9)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5669[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a7)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5645[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a6)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5633[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a4)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5609[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ab)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5693[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a1)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5573[13:0] );

									end
									else
									if((r_sys_run_step==9'h19b)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5477[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a5)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5621[13:0] );

									end
									else
									if((r_sys_run_step==9'h19c)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5489[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ae)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5729[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a8)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5657[13:0] );

									end
									else
									if((r_sys_run_step==9'h19d)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5525[13:0] );

									end
									else
									if((r_sys_run_step==9'h19e)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5537[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ad)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5717[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a3)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5597[13:0] );

									end
									else
									if((r_sys_run_step==9'h1af)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5741[13:0] );

									end
									else
									if((r_sys_run_step==9'h1aa)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5681[13:0] );

									end
									else
									if((r_sys_run_step==9'h1ac)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5705[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a0)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5561[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a2)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5585[13:0] );

									end
									else
									if((r_sys_run_step==9'h19f)) begin
										r_sub19_U_addr <= $signed( w_sys_tmp5549[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h19b<=r_sys_run_step && r_sys_run_step<=9'h1af)) begin
										r_sub19_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h19b<=r_sys_run_step && r_sys_run_step<=9'h1af)) begin
										r_sub19_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12867[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12857[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12862[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12897[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12907[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12932[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12872[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12937[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12882[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12902[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12927[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12912[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12942[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12917[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12887[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12947[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12877[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12922[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub19_result_addr <= $signed( w_sys_tmp12892[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub19_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h12)) begin
										r_sub19_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub19_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h9: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub09_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub09_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hda)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8746[13:0] );

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8656[13:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8668[13:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8704[13:0] );

									end
									else
									if((r_sys_run_step==9'hd9)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8740[13:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8710[13:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8752[13:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8680[13:0] );

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8650[13:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8662[13:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8716[13:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8620[13:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8722[13:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8692[13:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8728[13:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8626[13:0] );

									end
									else
									if((r_sys_run_step==9'hc9)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8644[13:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8674[13:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8698[13:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8686[13:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_sub09_T_addr <= $signed( w_sys_tmp8734[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hc7<=r_sys_run_step && r_sys_run_step<=9'hdb)) begin
										r_sub09_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hc7<=r_sys_run_step && r_sys_run_step<=9'hdb)) begin
										r_sub09_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc9)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp2981[13:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3065[13:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3029[13:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3017[13:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3077[13:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3089[13:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3041[13:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3161[13:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3125[13:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3053[13:0] );

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3005[13:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp2957[13:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp2969[13:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3113[13:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp2897[13:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp2909[13:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3101[13:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3149[13:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp2945[13:0] );

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp2993[13:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_sub09_V_addr <= $signed( w_sys_tmp3137[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hc4<=r_sys_run_step && r_sys_run_step<=9'hd8)) begin
										r_sub09_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hc4<=r_sys_run_step && r_sys_run_step<=9'hd8)) begin
										r_sub09_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc9)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp2981[13:0] );

									end
									else
									if((r_sys_run_step==9'hd0)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3065[13:0] );

									end
									else
									if((r_sys_run_step==9'hcd)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3029[13:0] );

									end
									else
									if((r_sys_run_step==9'hcc)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3017[13:0] );

									end
									else
									if((r_sys_run_step==9'hd1)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3077[13:0] );

									end
									else
									if((r_sys_run_step==9'hd2)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3089[13:0] );

									end
									else
									if((r_sys_run_step==9'hce)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3041[13:0] );

									end
									else
									if((r_sys_run_step==9'hd8)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3161[13:0] );

									end
									else
									if((r_sys_run_step==9'hd5)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3125[13:0] );

									end
									else
									if((r_sys_run_step==9'hcf)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3053[13:0] );

									end
									else
									if((r_sys_run_step==9'hcb)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3005[13:0] );

									end
									else
									if((r_sys_run_step==9'hc7)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp2957[13:0] );

									end
									else
									if((r_sys_run_step==9'hc8)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp2969[13:0] );

									end
									else
									if((r_sys_run_step==9'hd4)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3113[13:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp2897[13:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp2909[13:0] );

									end
									else
									if((r_sys_run_step==9'hd3)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3101[13:0] );

									end
									else
									if((r_sys_run_step==9'hd7)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3149[13:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp2945[13:0] );

									end
									else
									if((r_sys_run_step==9'hca)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp2993[13:0] );

									end
									else
									if((r_sys_run_step==9'hd6)) begin
										r_sub09_U_addr <= $signed( w_sys_tmp3137[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hc4<=r_sys_run_step && r_sys_run_step<=9'hd8)) begin
										r_sub09_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hc4<=r_sys_run_step && r_sys_run_step<=9'hd8)) begin
										r_sub09_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11912[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11957[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11882[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11887[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11892[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11927[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11942[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11932[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11867[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11872[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11937[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11922[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11907[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11877[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11947[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11917[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11952[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11902[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub09_result_addr <= $signed( w_sys_tmp11897[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub09_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h12)) begin
										r_sub09_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub09_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h8: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb8)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8542[13:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8548[13:0] );

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8602[13:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8572[13:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8494[13:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8512[13:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8488[13:0] );

									end
									else
									if((r_sys_run_step==9'hb4)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8518[13:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8566[13:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8530[13:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8524[13:0] );

									end
									else
									if((r_sys_run_step==9'hc4)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8614[13:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8578[13:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8608[13:0] );

									end
									else
									if((r_sys_run_step==9'hc5)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8620[13:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8596[13:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8554[13:0] );

									end
									else
									if((r_sys_run_step==9'hc6)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8626[13:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8590[13:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8560[13:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8536[13:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp8584[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hb1<=r_sys_run_step && r_sys_run_step<=9'hc6)) begin
										r_sub08_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hb1<=r_sys_run_step && r_sys_run_step<=9'hc6)) begin
										r_sub08_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb4)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2729[13:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2789[13:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2825[13:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2657[13:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2849[13:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2777[13:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2813[13:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2765[13:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2693[13:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2705[13:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2717[13:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2753[13:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2873[13:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2861[13:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2741[13:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2801[13:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2885[13:0] );

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2897[13:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2909[13:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2837[13:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp2681[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'haf<=r_sys_run_step && r_sys_run_step<=9'hc3)) begin
										r_sub08_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'haf<=r_sys_run_step && r_sys_run_step<=9'hc3)) begin
										r_sub08_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb4)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2729[13:0] );

									end
									else
									if((r_sys_run_step==9'hb9)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2789[13:0] );

									end
									else
									if((r_sys_run_step==9'hbc)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2825[13:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2657[13:0] );

									end
									else
									if((r_sys_run_step==9'hbe)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2849[13:0] );

									end
									else
									if((r_sys_run_step==9'hb8)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2777[13:0] );

									end
									else
									if((r_sys_run_step==9'hbb)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2813[13:0] );

									end
									else
									if((r_sys_run_step==9'hb7)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2765[13:0] );

									end
									else
									if((r_sys_run_step==9'hb1)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2693[13:0] );

									end
									else
									if((r_sys_run_step==9'hb2)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2705[13:0] );

									end
									else
									if((r_sys_run_step==9'hb3)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2717[13:0] );

									end
									else
									if((r_sys_run_step==9'hb6)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2753[13:0] );

									end
									else
									if((r_sys_run_step==9'hc0)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2873[13:0] );

									end
									else
									if((r_sys_run_step==9'hbf)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2861[13:0] );

									end
									else
									if((r_sys_run_step==9'hb5)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2741[13:0] );

									end
									else
									if((r_sys_run_step==9'hba)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2801[13:0] );

									end
									else
									if((r_sys_run_step==9'hc1)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2885[13:0] );

									end
									else
									if((r_sys_run_step==9'hc2)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2897[13:0] );

									end
									else
									if((r_sys_run_step==9'hc3)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2909[13:0] );

									end
									else
									if((r_sys_run_step==9'hbd)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2837[13:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp2681[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'haf<=r_sys_run_step && r_sys_run_step<=9'hc3)) begin
										r_sub08_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'haf<=r_sys_run_step && r_sys_run_step<=9'hc3)) begin
										r_sub08_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11782[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11812[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11832[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11842[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11777[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11797[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11767[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11772[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11822[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11802[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11827[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11792[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11807[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11862[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11857[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11787[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11852[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11847[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11817[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp11837[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h18: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub24_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub24_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5d)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10618[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10642[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10588[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10660[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10648[13:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10720[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10672[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10594[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10684[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10666[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10678[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10654[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10702[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10714[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10696[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10636[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10612[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10624[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10630[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10690[13:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_sub24_T_addr <= $signed( w_sys_tmp10708[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h5a<=r_sys_run_step && r_sys_run_step<=9'h6e)) begin
										r_sub24_T_datain <= w_sys_tmp10074;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h5a<=r_sys_run_step && r_sys_run_step<=9'h6e)) begin
										r_sub24_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h66)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6959[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6995[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp7019[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6923[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp7043[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp7007[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6911[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6791[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6983[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6887[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6899[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6827[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6863[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6875[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6971[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6935[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6839[13:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp7031[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6947[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6779[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_sub24_V_addr <= $signed( w_sys_tmp6851[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h59<=r_sys_run_step && r_sys_run_step<=9'h6d)) begin
										r_sub24_V_datain <= w_sys_tmp5767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h59<=r_sys_run_step && r_sys_run_step<=9'h6d)) begin
										r_sub24_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h66)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6959[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6995[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp7019[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6923[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp7043[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp7007[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6911[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6791[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6983[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6887[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6899[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6827[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6863[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6875[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6971[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6935[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6839[13:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp7031[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6947[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6779[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_sub24_U_addr <= $signed( w_sys_tmp6851[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h59<=r_sys_run_step && r_sys_run_step<=9'h6d)) begin
										r_sub24_U_datain <= w_sys_tmp5761;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h59<=r_sys_run_step && r_sys_run_step<=9'h6d)) begin
										r_sub24_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13468[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13383[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13438[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13403[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13418[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13423[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13458[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13408[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13413[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13433[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13448[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13443[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13378[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13388[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13393[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13428[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13398[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13463[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub24_result_addr <= $signed( w_sys_tmp13453[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub24_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h12)) begin
										r_sub24_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub24_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h16: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub22_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub22_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h38)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10396[13:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10450[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10426[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10390[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10384[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10324[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10378[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10402[13:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10456[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10372[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10414[13:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10444[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10360[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10462[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10408[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10330[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10432[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10366[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10348[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10438[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10420[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_sub22_T_addr <= $signed( w_sys_tmp10354[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2e<=r_sys_run_step && r_sys_run_step<=9'h43)) begin
										r_sub22_T_datain <= w_sys_tmp10074;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2e<=r_sys_run_step && r_sys_run_step<=9'h43)) begin
										r_sub22_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3a)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6431[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6323[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6479[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6383[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6371[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6419[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6311[13:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6515[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6491[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6347[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6335[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6263[13:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6527[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6395[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6455[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6359[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6443[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6407[13:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6503[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6251[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6299[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_sub22_V_addr <= $signed( w_sys_tmp6467[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2d<=r_sys_run_step && r_sys_run_step<=9'h42)) begin
										r_sub22_V_datain <= w_sys_tmp5767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2d<=r_sys_run_step && r_sys_run_step<=9'h42)) begin
										r_sub22_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3a)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6431[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6323[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6479[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6383[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6371[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6419[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6311[13:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6515[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6491[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6347[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6335[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6263[13:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6527[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6395[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6455[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6359[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6443[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6407[13:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6503[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6251[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6299[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_sub22_U_addr <= $signed( w_sys_tmp6467[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2d<=r_sys_run_step && r_sys_run_step<=9'h42)) begin
										r_sub22_U_datain <= w_sys_tmp5761;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2d<=r_sys_run_step && r_sys_run_step<=9'h42)) begin
										r_sub22_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13263[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13268[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13178[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13273[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13233[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13253[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13208[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13238[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13213[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13188[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13243[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13223[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13193[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13198[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13218[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13258[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13228[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13248[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13203[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub22_result_addr <= $signed( w_sys_tmp13183[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub22_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub22_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub22_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h17: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub23_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub23_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h58)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10588[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10558[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10522[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10570[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10486[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10504[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10528[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10510[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10594[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10492[13:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10582[13:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10576[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10546[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10456[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10498[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10540[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10564[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10552[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10462[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10516[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10534[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_sub23_T_addr <= $signed( w_sys_tmp10480[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h44<=r_sys_run_step && r_sys_run_step<=9'h59)) begin
										r_sub23_T_datain <= w_sys_tmp10074;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h44<=r_sys_run_step && r_sys_run_step<=9'h59)) begin
										r_sub23_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h53)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6731[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6743[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6575[13:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6767[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6755[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6683[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6659[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6515[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6587[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6635[13:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6791[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6599[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6611[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6527[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6671[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6695[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6563[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6647[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6707[13:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6779[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6719[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_sub23_V_addr <= $signed( w_sys_tmp6623[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h43<=r_sys_run_step && r_sys_run_step<=9'h58)) begin
										r_sub23_V_datain <= w_sys_tmp5767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h43<=r_sys_run_step && r_sys_run_step<=9'h58)) begin
										r_sub23_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h53)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6731[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6743[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6575[13:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6767[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6755[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6683[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6659[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6515[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6587[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6635[13:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6791[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6599[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6611[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6527[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6671[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6695[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6563[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6647[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6707[13:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6779[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6719[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_sub23_U_addr <= $signed( w_sys_tmp6623[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h43<=r_sys_run_step && r_sys_run_step<=9'h58)) begin
										r_sub23_U_datain <= w_sys_tmp5761;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h43<=r_sys_run_step && r_sys_run_step<=9'h58)) begin
										r_sub23_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13308[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13313[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13373[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13298[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13353[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13283[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13303[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13348[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13293[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13358[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13363[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13318[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13328[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13288[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13338[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13278[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13368[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13333[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13343[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub23_result_addr <= $signed( w_sys_tmp13323[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub23_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub23_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub23_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hc: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub12_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub12_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11c)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9142[13:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9016[13:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9088[13:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9106[13:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9034[13:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9052[13:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9136[13:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9046[13:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9010[13:0] );

									end
									else
									if((r_sys_run_step==9'h118)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9118[13:0] );

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9130[13:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9100[13:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9040[13:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9082[13:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9124[13:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9058[13:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9064[13:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9070[13:0] );

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9112[13:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9148[13:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9094[13:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_sub12_T_addr <= $signed( w_sys_tmp9076[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h108<=r_sys_run_step && r_sys_run_step<=9'h11d)) begin
										r_sub12_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h108<=r_sys_run_step && r_sys_run_step<=9'h11d)) begin
										r_sub12_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h118)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3929[13:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3797[13:0] );

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3917[13:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3905[13:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3857[13:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3677[13:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3737[13:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3809[13:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3833[13:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3821[13:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3749[13:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3665[13:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3773[13:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3941[13:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3785[13:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3881[13:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3761[13:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3713[13:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3893[13:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3869[13:0] );

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3725[13:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_sub12_V_addr <= $signed( w_sys_tmp3845[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h104<=r_sys_run_step && r_sys_run_step<=9'h119)) begin
										r_sub12_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h104<=r_sys_run_step && r_sys_run_step<=9'h119)) begin
										r_sub12_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h118)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3929[13:0] );

									end
									else
									if((r_sys_run_step==9'h10d)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3797[13:0] );

									end
									else
									if((r_sys_run_step==9'h117)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3917[13:0] );

									end
									else
									if((r_sys_run_step==9'h116)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3905[13:0] );

									end
									else
									if((r_sys_run_step==9'h112)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3857[13:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3677[13:0] );

									end
									else
									if((r_sys_run_step==9'h108)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3737[13:0] );

									end
									else
									if((r_sys_run_step==9'h10e)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3809[13:0] );

									end
									else
									if((r_sys_run_step==9'h110)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3833[13:0] );

									end
									else
									if((r_sys_run_step==9'h10f)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3821[13:0] );

									end
									else
									if((r_sys_run_step==9'h109)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3749[13:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3665[13:0] );

									end
									else
									if((r_sys_run_step==9'h10b)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3773[13:0] );

									end
									else
									if((r_sys_run_step==9'h119)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3941[13:0] );

									end
									else
									if((r_sys_run_step==9'h10c)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3785[13:0] );

									end
									else
									if((r_sys_run_step==9'h114)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3881[13:0] );

									end
									else
									if((r_sys_run_step==9'h10a)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3761[13:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3713[13:0] );

									end
									else
									if((r_sys_run_step==9'h115)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3893[13:0] );

									end
									else
									if((r_sys_run_step==9'h113)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3869[13:0] );

									end
									else
									if((r_sys_run_step==9'h107)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3725[13:0] );

									end
									else
									if((r_sys_run_step==9'h111)) begin
										r_sub12_U_addr <= $signed( w_sys_tmp3845[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h104<=r_sys_run_step && r_sys_run_step<=9'h119)) begin
										r_sub12_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h104<=r_sys_run_step && r_sys_run_step<=9'h119)) begin
										r_sub12_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12187[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12167[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12217[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12197[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12257[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12222[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12227[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12237[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12162[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12232[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12172[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12192[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12252[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12242[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12202[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12177[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12212[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12207[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12247[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub12_result_addr <= $signed( w_sys_tmp12182[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub12_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub12_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub12_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h3: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4f)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7912[13:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7954[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7918[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7936[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7942[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7858[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7972[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7834[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7840[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7864[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7924[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7948[13:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7960[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7930[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7906[13:0] );

									end
									else
									if((r_sys_run_step==9'h49)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7876[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7888[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7870[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7894[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7900[13:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7966[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp7882[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h44<=r_sys_run_step && r_sys_run_step<=9'h59)) begin
										r_sub03_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h44<=r_sys_run_step && r_sys_run_step<=9'h59)) begin
										r_sub03_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h49)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1445[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1457[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1505[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1469[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1541[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1529[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1409[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1421[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1361[13:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1601[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1433[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1565[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1385[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1481[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1517[13:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1625[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1553[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1397[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1493[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1589[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1577[13:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp1613[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h43<=r_sys_run_step && r_sys_run_step<=9'h58)) begin
										r_sub03_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h43<=r_sys_run_step && r_sys_run_step<=9'h58)) begin
										r_sub03_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h49)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1445[13:0] );

									end
									else
									if((r_sys_run_step==9'h4a)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1457[13:0] );

									end
									else
									if((r_sys_run_step==9'h4e)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1505[13:0] );

									end
									else
									if((r_sys_run_step==9'h4b)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1469[13:0] );

									end
									else
									if((r_sys_run_step==9'h51)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1541[13:0] );

									end
									else
									if((r_sys_run_step==9'h50)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1529[13:0] );

									end
									else
									if((r_sys_run_step==9'h46)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1409[13:0] );

									end
									else
									if((r_sys_run_step==9'h47)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1421[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1361[13:0] );

									end
									else
									if((r_sys_run_step==9'h56)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1601[13:0] );

									end
									else
									if((r_sys_run_step==9'h48)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1433[13:0] );

									end
									else
									if((r_sys_run_step==9'h53)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1565[13:0] );

									end
									else
									if((r_sys_run_step==9'h44)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1385[13:0] );

									end
									else
									if((r_sys_run_step==9'h4c)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1481[13:0] );

									end
									else
									if((r_sys_run_step==9'h4f)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1517[13:0] );

									end
									else
									if((r_sys_run_step==9'h58)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1625[13:0] );

									end
									else
									if((r_sys_run_step==9'h52)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1553[13:0] );

									end
									else
									if((r_sys_run_step==9'h45)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1397[13:0] );

									end
									else
									if((r_sys_run_step==9'h4d)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1493[13:0] );

									end
									else
									if((r_sys_run_step==9'h55)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1589[13:0] );

									end
									else
									if((r_sys_run_step==9'h54)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1577[13:0] );

									end
									else
									if((r_sys_run_step==9'h57)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp1613[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h43<=r_sys_run_step && r_sys_run_step<=9'h58)) begin
										r_sub03_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h43<=r_sys_run_step && r_sys_run_step<=9'h58)) begin
										r_sub03_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11352[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11267[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11297[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11322[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11302[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11342[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11337[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11307[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11347[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11287[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11332[13:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11362[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11282[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11292[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11277[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11257[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11312[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11317[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11357[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11272[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp11327[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h14)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h2: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3e)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7810[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7792[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7756[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7732[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7816[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7786[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7738[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7750[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7744[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7768[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7702[13:0] );

									end
									else
									if((r_sys_run_step==9'h43)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7840[13:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7834[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7804[13:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7822[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7774[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7726[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7780[13:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7828[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7798[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7708[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp7762[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2e<=r_sys_run_step && r_sys_run_step<=9'h43)) begin
										r_sub02_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2e<=r_sys_run_step && r_sys_run_step<=9'h43)) begin
										r_sub02_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2e)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1097[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1229[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1313[13:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1361[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1289[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1277[13:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1349[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1253[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1193[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1241[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1181[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1205[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1265[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1145[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1169[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1217[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1301[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1109[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1157[13:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1337[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp1325[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2e<=r_sys_run_step && r_sys_run_step<=9'h42)) begin
										r_sub02_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2e<=r_sys_run_step && r_sys_run_step<=9'h42)) begin
										r_sub02_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2e)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1097[13:0] );

									end
									else
									if((r_sys_run_step==9'h37)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1229[13:0] );

									end
									else
									if((r_sys_run_step==9'h3e)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1313[13:0] );

									end
									else
									if((r_sys_run_step==9'h42)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1361[13:0] );

									end
									else
									if((r_sys_run_step==9'h3c)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1289[13:0] );

									end
									else
									if((r_sys_run_step==9'h3b)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1277[13:0] );

									end
									else
									if((r_sys_run_step==9'h41)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1349[13:0] );

									end
									else
									if((r_sys_run_step==9'h39)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1253[13:0] );

									end
									else
									if((r_sys_run_step==9'h34)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1193[13:0] );

									end
									else
									if((r_sys_run_step==9'h38)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1241[13:0] );

									end
									else
									if((r_sys_run_step==9'h33)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1181[13:0] );

									end
									else
									if((r_sys_run_step==9'h35)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1205[13:0] );

									end
									else
									if((r_sys_run_step==9'h3a)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1265[13:0] );

									end
									else
									if((r_sys_run_step==9'h30)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1145[13:0] );

									end
									else
									if((r_sys_run_step==9'h32)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1169[13:0] );

									end
									else
									if((r_sys_run_step==9'h36)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1217[13:0] );

									end
									else
									if((r_sys_run_step==9'h3d)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1301[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1109[13:0] );

									end
									else
									if((r_sys_run_step==9'h31)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1157[13:0] );

									end
									else
									if((r_sys_run_step==9'h40)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1337[13:0] );

									end
									else
									if((r_sys_run_step==9'h3f)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp1325[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2e<=r_sys_run_step && r_sys_run_step<=9'h42)) begin
										r_sub02_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2e<=r_sys_run_step && r_sys_run_step<=9'h42)) begin
										r_sub02_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11007[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11182[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10840[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11237[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10972[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10846[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10952[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10927[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10967[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11177[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10828[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11217[13:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10987[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11167[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10810[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10804[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10957[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11172[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10937[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10932[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10977[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10962[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11012[13:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10997[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11207[13:0] );

									end
									else
									if((r_sys_run_step==9'h2e)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11252[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11192[13:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11242[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11222[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11227[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11017[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11232[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10822[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11202[13:0] );

									end
									else
									if((r_sys_run_step==9'h2f)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11257[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11212[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10834[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10947[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11247[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10942[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11162[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11197[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11002[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10922[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10816[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp11187[13:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10982[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp10992[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h2f)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hb: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub11_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub11_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h107)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp9016[13:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8956[13:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8878[13:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8908[13:0] );

									end
									else
									if((r_sys_run_step==9'h104)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8998[13:0] );

									end
									else
									if((r_sys_run_step==9'h105)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp9004[13:0] );

									end
									else
									if((r_sys_run_step==9'hf6)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8914[13:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8980[13:0] );

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8974[13:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8884[13:0] );

									end
									else
									if((r_sys_run_step==9'h106)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp9010[13:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8938[13:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8944[13:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8968[13:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8926[13:0] );

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8992[13:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8902[13:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8950[13:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8962[13:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8920[13:0] );

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8986[13:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_sub11_T_addr <= $signed( w_sys_tmp8932[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hf2<=r_sys_run_step && r_sys_run_step<=9'h107)) begin
										r_sub11_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hf2<=r_sys_run_step && r_sys_run_step<=9'h107)) begin
										r_sub11_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf6)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3521[13:0] );

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3641[13:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3653[13:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3461[13:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3413[13:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3509[13:0] );

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3677[13:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3497[13:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3617[13:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3473[13:0] );

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3665[13:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3533[13:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3581[13:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3569[13:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3557[13:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3629[13:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3593[13:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3485[13:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3437[13:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3545[13:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3449[13:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_sub11_V_addr <= $signed( w_sys_tmp3605[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hee<=r_sys_run_step && r_sys_run_step<=9'h103)) begin
										r_sub11_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hee<=r_sys_run_step && r_sys_run_step<=9'h103)) begin
										r_sub11_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf6)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3521[13:0] );

									end
									else
									if((r_sys_run_step==9'h100)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3641[13:0] );

									end
									else
									if((r_sys_run_step==9'h101)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3653[13:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3461[13:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3413[13:0] );

									end
									else
									if((r_sys_run_step==9'hf5)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3509[13:0] );

									end
									else
									if((r_sys_run_step==9'h103)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3677[13:0] );

									end
									else
									if((r_sys_run_step==9'hf4)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3497[13:0] );

									end
									else
									if((r_sys_run_step==9'hfe)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3617[13:0] );

									end
									else
									if((r_sys_run_step==9'hf2)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3473[13:0] );

									end
									else
									if((r_sys_run_step==9'h102)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3665[13:0] );

									end
									else
									if((r_sys_run_step==9'hf7)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3533[13:0] );

									end
									else
									if((r_sys_run_step==9'hfb)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3581[13:0] );

									end
									else
									if((r_sys_run_step==9'hfa)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3569[13:0] );

									end
									else
									if((r_sys_run_step==9'hf9)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3557[13:0] );

									end
									else
									if((r_sys_run_step==9'hff)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3629[13:0] );

									end
									else
									if((r_sys_run_step==9'hfc)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3593[13:0] );

									end
									else
									if((r_sys_run_step==9'hf3)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3485[13:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3437[13:0] );

									end
									else
									if((r_sys_run_step==9'hf8)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3545[13:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3449[13:0] );

									end
									else
									if((r_sys_run_step==9'hfd)) begin
										r_sub11_U_addr <= $signed( w_sys_tmp3605[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hee<=r_sys_run_step && r_sys_run_step<=9'h103)) begin
										r_sub11_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hee<=r_sys_run_step && r_sys_run_step<=9'h103)) begin
										r_sub11_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12097[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12087[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12117[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12077[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12157[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12102[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12112[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12132[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12062[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12147[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12067[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12127[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12082[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12107[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12152[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12142[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12122[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12092[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12137[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub11_result_addr <= $signed( w_sys_tmp12072[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub11_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub11_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub11_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'he: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub14_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub14_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h144)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9382[13:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9364[13:0] );

									end
									else
									if((r_sys_run_step==9'h13b)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9328[13:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9388[13:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9316[13:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9334[13:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9274[13:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9280[13:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9370[13:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9340[13:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9304[13:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9358[13:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9346[13:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9406[13:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9322[13:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9298[13:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9310[13:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9394[13:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9376[13:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9400[13:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_sub14_T_addr <= $signed( w_sys_tmp9352[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h134<=r_sys_run_step && r_sys_run_step<=9'h148)) begin
										r_sub14_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h134<=r_sys_run_step && r_sys_run_step<=9'h148)) begin
										r_sub14_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13b)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4349[13:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4385[13:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4433[13:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4325[13:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4409[13:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4373[13:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4337[13:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4301[13:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4421[13:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4277[13:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4361[13:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4445[13:0] );

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4181[13:0] );

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4193[13:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4289[13:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4229[13:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4241[13:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4397[13:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4253[13:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4265[13:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_sub14_V_addr <= $signed( w_sys_tmp4313[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h12f<=r_sys_run_step && r_sys_run_step<=9'h143)) begin
										r_sub14_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h12f<=r_sys_run_step && r_sys_run_step<=9'h143)) begin
										r_sub14_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13b)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4349[13:0] );

									end
									else
									if((r_sys_run_step==9'h13e)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4385[13:0] );

									end
									else
									if((r_sys_run_step==9'h142)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4433[13:0] );

									end
									else
									if((r_sys_run_step==9'h139)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4325[13:0] );

									end
									else
									if((r_sys_run_step==9'h140)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4409[13:0] );

									end
									else
									if((r_sys_run_step==9'h13d)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4373[13:0] );

									end
									else
									if((r_sys_run_step==9'h13a)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4337[13:0] );

									end
									else
									if((r_sys_run_step==9'h137)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4301[13:0] );

									end
									else
									if((r_sys_run_step==9'h141)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4421[13:0] );

									end
									else
									if((r_sys_run_step==9'h135)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4277[13:0] );

									end
									else
									if((r_sys_run_step==9'h13c)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4361[13:0] );

									end
									else
									if((r_sys_run_step==9'h143)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4445[13:0] );

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4181[13:0] );

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4193[13:0] );

									end
									else
									if((r_sys_run_step==9'h136)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4289[13:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4229[13:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4241[13:0] );

									end
									else
									if((r_sys_run_step==9'h13f)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4397[13:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4253[13:0] );

									end
									else
									if((r_sys_run_step==9'h134)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4265[13:0] );

									end
									else
									if((r_sys_run_step==9'h138)) begin
										r_sub14_U_addr <= $signed( w_sys_tmp4313[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h12f<=r_sys_run_step && r_sys_run_step<=9'h143)) begin
										r_sub14_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h12f<=r_sys_run_step && r_sys_run_step<=9'h143)) begin
										r_sub14_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12372[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12382[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12407[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12432[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12447[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12367[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12442[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12377[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12412[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12402[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12392[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12452[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12422[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12387[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12437[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12397[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12362[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12417[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub14_result_addr <= $signed( w_sys_tmp12427[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub14_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h12)) begin
										r_sub14_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub14_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h1: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2a)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7690[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7570[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7666[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7612[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7642[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7618[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7600[13:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7702[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7678[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7696[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7594[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7576[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7660[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7624[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7630[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7654[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7672[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7708[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7684[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7606[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7636[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp7648[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h18<=r_sys_run_step && r_sys_run_step<=9'h2d)) begin
										r_sub01_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h18<=r_sys_run_step && r_sys_run_step<=9'h2d)) begin
										r_sub01_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h28)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp1049[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp917[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp941[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp1061[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp953[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp1013[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp1025[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp989[13:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp1097[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp965[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp1073[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp881[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp893[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp833[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp929[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp905[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp977[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp845[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp1001[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp1085[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp1109[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp1037[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h18<=r_sys_run_step && r_sys_run_step<=9'h2d)) begin
										r_sub01_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h18<=r_sys_run_step && r_sys_run_step<=9'h2d)) begin
										r_sub01_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h28)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp1049[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp917[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp941[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp1061[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp953[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp1013[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp1025[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp989[13:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp1097[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp965[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp1073[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp881[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp893[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp833[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp929[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp905[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp977[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp845[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp1001[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp1085[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp1109[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp1037[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h18<=r_sys_run_step && r_sys_run_step<=9'h2d)) begin
										r_sub01_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h18<=r_sys_run_step && r_sys_run_step<=9'h2d)) begin
										r_sub01_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp11007[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10840[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10972[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10780[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10846[13:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10952[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10768[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10927[13:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10967[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10828[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10987[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10798[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10810[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10804[13:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10957[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10932[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10937[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10977[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10774[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10962[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp11012[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10997[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10786[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp11017[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10792[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10822[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10834[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10947[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10942[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp11002[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10816[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10922[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10992[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp10982[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h21)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7534[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7468[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7570[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7456[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7522[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7462[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7486[13:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7576[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7552[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7492[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7546[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7504[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7450[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7510[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7474[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7540[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7480[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7516[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7528[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7498[13:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7564[13:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp7558[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h17)) begin
										r_sub00_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h17)) begin
										r_sub00_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp641[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp797[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp593[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp689[13:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp809[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp725[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp761[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp749[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp605[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp833[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp617[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp653[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp629[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp665[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp785[13:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp845[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp773[13:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp821[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp737[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp677[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp701[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp713[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h17)) begin
										r_sub00_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h17)) begin
										r_sub00_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp641[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp797[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp593[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp689[13:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp809[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp725[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp761[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp749[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp605[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp833[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp617[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp653[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp629[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp665[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp785[13:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp845[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp773[13:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp821[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp737[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp677[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp701[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp713[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h17)) begin
										r_sub00_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h17)) begin
										r_sub00_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10738[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10774[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10756[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10840[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10786[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10780[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10762[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10792[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10846[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10822[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10744[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10768[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10834[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10750[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10828[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10798[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10816[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10810[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10804[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp10732[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hd: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub13_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub13_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11e)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9142[13:0] );

									end
									else
									if((r_sys_run_step==9'h130)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9262[13:0] );

									end
									else
									if((r_sys_run_step==9'h12e)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9250[13:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9226[13:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9172[13:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9220[13:0] );

									end
									else
									if((r_sys_run_step==9'h133)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9280[13:0] );

									end
									else
									if((r_sys_run_step==9'h132)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9274[13:0] );

									end
									else
									if((r_sys_run_step==9'h131)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9268[13:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9214[13:0] );

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9238[13:0] );

									end
									else
									if((r_sys_run_step==9'h12d)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9244[13:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9196[13:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9208[13:0] );

									end
									else
									if((r_sys_run_step==9'h12f)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9256[13:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9184[13:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9166[13:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9178[13:0] );

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9232[13:0] );

									end
									else
									if((r_sys_run_step==9'h124)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9190[13:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9202[13:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_sub13_T_addr <= $signed( w_sys_tmp9148[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h11e<=r_sys_run_step && r_sys_run_step<=9'h133)) begin
										r_sub13_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h11e<=r_sys_run_step && r_sys_run_step<=9'h133)) begin
										r_sub13_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h124)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4073[13:0] );

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4157[13:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4049[13:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4025[13:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4097[13:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4061[13:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4145[13:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4001[13:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp3989[13:0] );

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4169[13:0] );

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp3941[13:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp3965[13:0] );

									end
									else
									if((r_sys_run_step==9'h12e)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4193[13:0] );

									end
									else
									if((r_sys_run_step==9'h12d)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4181[13:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4037[13:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4133[13:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4121[13:0] );

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp3977[13:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4013[13:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4085[13:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_sub13_V_addr <= $signed( w_sys_tmp4109[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h11a<=r_sys_run_step && r_sys_run_step<=9'h12e)) begin
										r_sub13_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h11a<=r_sys_run_step && r_sys_run_step<=9'h12e)) begin
										r_sub13_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h124)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4073[13:0] );

									end
									else
									if((r_sys_run_step==9'h12b)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4157[13:0] );

									end
									else
									if((r_sys_run_step==9'h122)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4049[13:0] );

									end
									else
									if((r_sys_run_step==9'h120)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4025[13:0] );

									end
									else
									if((r_sys_run_step==9'h126)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4097[13:0] );

									end
									else
									if((r_sys_run_step==9'h123)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4061[13:0] );

									end
									else
									if((r_sys_run_step==9'h12a)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4145[13:0] );

									end
									else
									if((r_sys_run_step==9'h11e)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4001[13:0] );

									end
									else
									if((r_sys_run_step==9'h11d)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp3989[13:0] );

									end
									else
									if((r_sys_run_step==9'h12c)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4169[13:0] );

									end
									else
									if((r_sys_run_step==9'h11a)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp3941[13:0] );

									end
									else
									if((r_sys_run_step==9'h11b)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp3965[13:0] );

									end
									else
									if((r_sys_run_step==9'h12e)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4193[13:0] );

									end
									else
									if((r_sys_run_step==9'h12d)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4181[13:0] );

									end
									else
									if((r_sys_run_step==9'h121)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4037[13:0] );

									end
									else
									if((r_sys_run_step==9'h129)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4133[13:0] );

									end
									else
									if((r_sys_run_step==9'h128)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4121[13:0] );

									end
									else
									if((r_sys_run_step==9'h11c)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp3977[13:0] );

									end
									else
									if((r_sys_run_step==9'h11f)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4013[13:0] );

									end
									else
									if((r_sys_run_step==9'h125)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4085[13:0] );

									end
									else
									if((r_sys_run_step==9'h127)) begin
										r_sub13_U_addr <= $signed( w_sys_tmp4109[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h11a<=r_sys_run_step && r_sys_run_step<=9'h12e)) begin
										r_sub13_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h11a<=r_sys_run_step && r_sys_run_step<=9'h12e)) begin
										r_sub13_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12342[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12262[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12292[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12282[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12287[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12347[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12272[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12352[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12297[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12267[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12322[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12277[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12302[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12317[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12337[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12327[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12357[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12332[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12307[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub13_result_addr <= $signed( w_sys_tmp12312[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub13_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub13_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub13_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h7: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9d)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8380[13:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8458[13:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8356[13:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8470[13:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8446[13:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8392[13:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8398[13:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8428[13:0] );

									end
									else
									if((r_sys_run_step==9'hb0)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8494[13:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8452[13:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8362[13:0] );

									end
									else
									if((r_sys_run_step==9'haf)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8488[13:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8440[13:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8482[13:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8422[13:0] );

									end
									else
									if((r_sys_run_step==9'ha6)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8434[13:0] );

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8476[13:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8464[13:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8416[13:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8404[13:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8386[13:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp8410[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h9b<=r_sys_run_step && r_sys_run_step<=9'hb0)) begin
										r_sub07_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h9b<=r_sys_run_step && r_sys_run_step<=9'hb0)) begin
										r_sub07_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha6)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2561[13:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2549[13:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2393[13:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2381[13:0] );

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2645[13:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2597[13:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2621[13:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2573[13:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2525[13:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2441[13:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2657[13:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2609[13:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2501[13:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2465[13:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2489[13:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2585[13:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2513[13:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2453[13:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2429[13:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2477[13:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2537[13:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp2633[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h99<=r_sys_run_step && r_sys_run_step<=9'hae)) begin
										r_sub07_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h99<=r_sys_run_step && r_sys_run_step<=9'hae)) begin
										r_sub07_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha6)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2561[13:0] );

									end
									else
									if((r_sys_run_step==9'ha5)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2549[13:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2393[13:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2381[13:0] );

									end
									else
									if((r_sys_run_step==9'had)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2645[13:0] );

									end
									else
									if((r_sys_run_step==9'ha9)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2597[13:0] );

									end
									else
									if((r_sys_run_step==9'hab)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2621[13:0] );

									end
									else
									if((r_sys_run_step==9'ha7)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2573[13:0] );

									end
									else
									if((r_sys_run_step==9'ha3)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2525[13:0] );

									end
									else
									if((r_sys_run_step==9'h9c)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2441[13:0] );

									end
									else
									if((r_sys_run_step==9'hae)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2657[13:0] );

									end
									else
									if((r_sys_run_step==9'haa)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2609[13:0] );

									end
									else
									if((r_sys_run_step==9'ha1)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2501[13:0] );

									end
									else
									if((r_sys_run_step==9'h9e)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2465[13:0] );

									end
									else
									if((r_sys_run_step==9'ha0)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2489[13:0] );

									end
									else
									if((r_sys_run_step==9'ha8)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2585[13:0] );

									end
									else
									if((r_sys_run_step==9'ha2)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2513[13:0] );

									end
									else
									if((r_sys_run_step==9'h9d)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2453[13:0] );

									end
									else
									if((r_sys_run_step==9'h9b)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2429[13:0] );

									end
									else
									if((r_sys_run_step==9'h9f)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2477[13:0] );

									end
									else
									if((r_sys_run_step==9'ha4)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2537[13:0] );

									end
									else
									if((r_sys_run_step==9'hac)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp2633[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h99<=r_sys_run_step && r_sys_run_step<=9'hae)) begin
										r_sub07_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h99<=r_sys_run_step && r_sys_run_step<=9'hae)) begin
										r_sub07_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11762[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11682[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11677[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11717[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11737[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11702[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11757[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11752[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11667[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11672[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11742[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11692[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11697[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11727[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11712[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11747[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11732[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11722[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11687[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp11707[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h10: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub16_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub16_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h162)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9562[13:0] );

									end
									else
									if((r_sys_run_step==9'h161)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9556[13:0] );

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9670[13:0] );

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9634[13:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9610[13:0] );

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9664[13:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9598[13:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9646[13:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9574[13:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9604[13:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9532[13:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9640[13:0] );

									end
									else
									if((r_sys_run_step==9'h172)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9658[13:0] );

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9628[13:0] );

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9622[13:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9580[13:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9568[13:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9538[13:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9592[13:0] );

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9616[13:0] );

									end
									else
									if((r_sys_run_step==9'h171)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9652[13:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_sub16_T_addr <= $signed( w_sys_tmp9586[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h15f<=r_sys_run_step && r_sys_run_step<=9'h174)) begin
										r_sub16_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h15f<=r_sys_run_step && r_sys_run_step<=9'h174)) begin
										r_sub16_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h161)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4805[13:0] );

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4949[13:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4913[13:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4721[13:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4829[13:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4889[13:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4877[13:0] );

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4925[13:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4853[13:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4901[13:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4865[13:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4817[13:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4841[13:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4757[13:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4745[13:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4769[13:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4697[13:0] );

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4937[13:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4733[13:0] );

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4961[13:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4781[13:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_sub16_V_addr <= $signed( w_sys_tmp4793[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h159<=r_sys_run_step && r_sys_run_step<=9'h16e)) begin
										r_sub16_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h159<=r_sys_run_step && r_sys_run_step<=9'h16e)) begin
										r_sub16_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h161)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4805[13:0] );

									end
									else
									if((r_sys_run_step==9'h16d)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4949[13:0] );

									end
									else
									if((r_sys_run_step==9'h16a)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4913[13:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4721[13:0] );

									end
									else
									if((r_sys_run_step==9'h163)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4829[13:0] );

									end
									else
									if((r_sys_run_step==9'h168)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4889[13:0] );

									end
									else
									if((r_sys_run_step==9'h167)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4877[13:0] );

									end
									else
									if((r_sys_run_step==9'h16b)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4925[13:0] );

									end
									else
									if((r_sys_run_step==9'h165)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4853[13:0] );

									end
									else
									if((r_sys_run_step==9'h169)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4901[13:0] );

									end
									else
									if((r_sys_run_step==9'h166)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4865[13:0] );

									end
									else
									if((r_sys_run_step==9'h162)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4817[13:0] );

									end
									else
									if((r_sys_run_step==9'h164)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4841[13:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4757[13:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4745[13:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4769[13:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4697[13:0] );

									end
									else
									if((r_sys_run_step==9'h16c)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4937[13:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4733[13:0] );

									end
									else
									if((r_sys_run_step==9'h16e)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4961[13:0] );

									end
									else
									if((r_sys_run_step==9'h15f)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4781[13:0] );

									end
									else
									if((r_sys_run_step==9'h160)) begin
										r_sub16_U_addr <= $signed( w_sys_tmp4793[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h159<=r_sys_run_step && r_sys_run_step<=9'h16e)) begin
										r_sub16_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h159<=r_sys_run_step && r_sys_run_step<=9'h16e)) begin
										r_sub16_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12592[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12572[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12647[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12607[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12652[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12567[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12612[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12597[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12622[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12617[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12577[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12602[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12627[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12632[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12557[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12582[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12587[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12642[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12562[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub16_result_addr <= $signed( w_sys_tmp12637[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub16_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub16_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub16_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h6: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h98)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8350[13:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8284[13:0] );

									end
									else
									if((r_sys_run_step==9'h99)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8356[13:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8320[13:0] );

									end
									else
									if((r_sys_run_step==9'h85)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8224[13:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8332[13:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8260[13:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8248[13:0] );

									end
									else
									if((r_sys_run_step==9'h9a)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8362[13:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8254[13:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8290[13:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8278[13:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8302[13:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8338[13:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8272[13:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8266[13:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8230[13:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8296[13:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8326[13:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8308[13:0] );

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8344[13:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp8314[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h85<=r_sys_run_step && r_sys_run_step<=9'h9a)) begin
										r_sub06_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h85<=r_sys_run_step && r_sys_run_step<=9'h9a)) begin
										r_sub06_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h85)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2165[13:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2273[13:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2285[13:0] );

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2393[13:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2261[13:0] );

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2381[13:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2177[13:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2189[13:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2213[13:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2129[13:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2249[13:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2369[13:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2333[13:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2225[13:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2201[13:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2357[13:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2237[13:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2321[13:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2309[13:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2345[13:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2153[13:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp2297[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h83<=r_sys_run_step && r_sys_run_step<=9'h98)) begin
										r_sub06_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h83<=r_sys_run_step && r_sys_run_step<=9'h98)) begin
										r_sub06_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h85)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2165[13:0] );

									end
									else
									if((r_sys_run_step==9'h8e)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2273[13:0] );

									end
									else
									if((r_sys_run_step==9'h8f)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2285[13:0] );

									end
									else
									if((r_sys_run_step==9'h98)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2393[13:0] );

									end
									else
									if((r_sys_run_step==9'h8d)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2261[13:0] );

									end
									else
									if((r_sys_run_step==9'h97)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2381[13:0] );

									end
									else
									if((r_sys_run_step==9'h86)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2177[13:0] );

									end
									else
									if((r_sys_run_step==9'h87)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2189[13:0] );

									end
									else
									if((r_sys_run_step==9'h89)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2213[13:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2129[13:0] );

									end
									else
									if((r_sys_run_step==9'h8c)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2249[13:0] );

									end
									else
									if((r_sys_run_step==9'h96)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2369[13:0] );

									end
									else
									if((r_sys_run_step==9'h93)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2333[13:0] );

									end
									else
									if((r_sys_run_step==9'h8a)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2225[13:0] );

									end
									else
									if((r_sys_run_step==9'h88)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2201[13:0] );

									end
									else
									if((r_sys_run_step==9'h95)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2357[13:0] );

									end
									else
									if((r_sys_run_step==9'h8b)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2237[13:0] );

									end
									else
									if((r_sys_run_step==9'h92)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2321[13:0] );

									end
									else
									if((r_sys_run_step==9'h91)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2309[13:0] );

									end
									else
									if((r_sys_run_step==9'h94)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2345[13:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2153[13:0] );

									end
									else
									if((r_sys_run_step==9'h90)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp2297[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h83<=r_sys_run_step && r_sys_run_step<=9'h98)) begin
										r_sub06_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h83<=r_sys_run_step && r_sys_run_step<=9'h98)) begin
										r_sub06_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11572[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11652[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11627[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11602[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11647[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11597[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11642[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11607[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11622[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11612[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11662[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11657[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11567[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11617[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11592[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11582[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11632[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11587[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11577[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp11637[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'hf: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub15_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub15_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h155)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9484[13:0] );

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9490[13:0] );

									end
									else
									if((r_sys_run_step==9'h15c)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9526[13:0] );

									end
									else
									if((r_sys_run_step==9'h15b)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9520[13:0] );

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9460[13:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9472[13:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9436[13:0] );

									end
									else
									if((r_sys_run_step==9'h157)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9496[13:0] );

									end
									else
									if((r_sys_run_step==9'h15a)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9514[13:0] );

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9466[13:0] );

									end
									else
									if((r_sys_run_step==9'h15d)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9532[13:0] );

									end
									else
									if((r_sys_run_step==9'h159)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9508[13:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9424[13:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9478[13:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9502[13:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9430[13:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9442[13:0] );

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9448[13:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9418[13:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9412[13:0] );

									end
									else
									if((r_sys_run_step==9'h15e)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9538[13:0] );

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_sub15_T_addr <= $signed( w_sys_tmp9454[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h149<=r_sys_run_step && r_sys_run_step<=9'h15e)) begin
										r_sub15_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h149<=r_sys_run_step && r_sys_run_step<=9'h15e)) begin
										r_sub15_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h157)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4685[13:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4481[13:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4457[13:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4505[13:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4565[13:0] );

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4589[13:0] );

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4601[13:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4493[13:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4529[13:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4577[13:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4517[13:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4553[13:0] );

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4625[13:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4649[13:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4541[13:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4697[13:0] );

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4613[13:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4637[13:0] );

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4673[13:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4661[13:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_sub15_V_addr <= $signed( w_sys_tmp4469[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h144<=r_sys_run_step && r_sys_run_step<=9'h158)) begin
										r_sub15_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h144<=r_sys_run_step && r_sys_run_step<=9'h158)) begin
										r_sub15_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h157)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4685[13:0] );

									end
									else
									if((r_sys_run_step==9'h146)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4481[13:0] );

									end
									else
									if((r_sys_run_step==9'h144)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4457[13:0] );

									end
									else
									if((r_sys_run_step==9'h148)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4505[13:0] );

									end
									else
									if((r_sys_run_step==9'h14d)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4565[13:0] );

									end
									else
									if((r_sys_run_step==9'h14f)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4589[13:0] );

									end
									else
									if((r_sys_run_step==9'h150)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4601[13:0] );

									end
									else
									if((r_sys_run_step==9'h147)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4493[13:0] );

									end
									else
									if((r_sys_run_step==9'h14a)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4529[13:0] );

									end
									else
									if((r_sys_run_step==9'h14e)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4577[13:0] );

									end
									else
									if((r_sys_run_step==9'h149)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4517[13:0] );

									end
									else
									if((r_sys_run_step==9'h14c)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4553[13:0] );

									end
									else
									if((r_sys_run_step==9'h152)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4625[13:0] );

									end
									else
									if((r_sys_run_step==9'h154)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4649[13:0] );

									end
									else
									if((r_sys_run_step==9'h14b)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4541[13:0] );

									end
									else
									if((r_sys_run_step==9'h158)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4697[13:0] );

									end
									else
									if((r_sys_run_step==9'h151)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4613[13:0] );

									end
									else
									if((r_sys_run_step==9'h153)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4637[13:0] );

									end
									else
									if((r_sys_run_step==9'h156)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4673[13:0] );

									end
									else
									if((r_sys_run_step==9'h155)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4661[13:0] );

									end
									else
									if((r_sys_run_step==9'h145)) begin
										r_sub15_U_addr <= $signed( w_sys_tmp4469[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h144<=r_sys_run_step && r_sys_run_step<=9'h158)) begin
										r_sub15_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h144<=r_sys_run_step && r_sys_run_step<=9'h158)) begin
										r_sub15_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12457[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12502[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12547[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12532[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12507[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12517[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12482[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12497[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12462[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12487[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12522[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12537[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12512[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12527[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12467[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12472[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12477[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12542[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12492[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub15_result_addr <= $signed( w_sys_tmp12552[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub15_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub15_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub15_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h5: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7e)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8194[13:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8104[13:0] );

									end
									else
									if((r_sys_run_step==9'h83)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8224[13:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8146[13:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8128[13:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8164[13:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8116[13:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8170[13:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8200[13:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8110[13:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8206[13:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8134[13:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8152[13:0] );

									end
									else
									if((r_sys_run_step==9'h7b)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8176[13:0] );

									end
									else
									if((r_sys_run_step==9'h84)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8230[13:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8188[13:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8218[13:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8212[13:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8122[13:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8158[13:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8182[13:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp8140[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h6f<=r_sys_run_step && r_sys_run_step<=9'h84)) begin
										r_sub05_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h6f<=r_sys_run_step && r_sys_run_step<=9'h84)) begin
										r_sub05_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7b)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2045[13:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2069[13:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1961[13:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1889[13:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2033[13:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1925[13:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1937[13:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2021[13:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2129[13:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1997[13:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2105[13:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2009[13:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1901[13:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2081[13:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2117[13:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1985[13:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1949[13:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1973[13:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2093[13:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp2057[13:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1913[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h6e<=r_sys_run_step && r_sys_run_step<=9'h82)) begin
										r_sub05_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h6e<=r_sys_run_step && r_sys_run_step<=9'h82)) begin
										r_sub05_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7b)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2045[13:0] );

									end
									else
									if((r_sys_run_step==9'h7d)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2069[13:0] );

									end
									else
									if((r_sys_run_step==9'h74)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1961[13:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1889[13:0] );

									end
									else
									if((r_sys_run_step==9'h7a)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2033[13:0] );

									end
									else
									if((r_sys_run_step==9'h71)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1925[13:0] );

									end
									else
									if((r_sys_run_step==9'h72)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1937[13:0] );

									end
									else
									if((r_sys_run_step==9'h79)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2021[13:0] );

									end
									else
									if((r_sys_run_step==9'h82)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2129[13:0] );

									end
									else
									if((r_sys_run_step==9'h77)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1997[13:0] );

									end
									else
									if((r_sys_run_step==9'h80)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2105[13:0] );

									end
									else
									if((r_sys_run_step==9'h78)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2009[13:0] );

									end
									else
									if((r_sys_run_step==9'h6f)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1901[13:0] );

									end
									else
									if((r_sys_run_step==9'h7e)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2081[13:0] );

									end
									else
									if((r_sys_run_step==9'h81)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2117[13:0] );

									end
									else
									if((r_sys_run_step==9'h76)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1985[13:0] );

									end
									else
									if((r_sys_run_step==9'h73)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1949[13:0] );

									end
									else
									if((r_sys_run_step==9'h75)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1973[13:0] );

									end
									else
									if((r_sys_run_step==9'h7f)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2093[13:0] );

									end
									else
									if((r_sys_run_step==9'h7c)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp2057[13:0] );

									end
									else
									if((r_sys_run_step==9'h70)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1913[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h6e<=r_sys_run_step && r_sys_run_step<=9'h82)) begin
										r_sub05_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h6e<=r_sys_run_step && r_sys_run_step<=9'h82)) begin
										r_sub05_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11512[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11522[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11472[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11482[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11552[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11562[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11487[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11467[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11492[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11557[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11507[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11537[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11477[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11542[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11527[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11532[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11497[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11547[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11502[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp11517[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h12: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub18_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub18_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h191)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9844[13:0] );

									end
									else
									if((r_sys_run_step==9'h19f)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9928[13:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9856[13:0] );

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9862[13:0] );

									end
									else
									if((r_sys_run_step==9'h19d)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9916[13:0] );

									end
									else
									if((r_sys_run_step==9'h19c)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9910[13:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9796[13:0] );

									end
									else
									if((r_sys_run_step==9'h19a)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9898[13:0] );

									end
									else
									if((r_sys_run_step==9'h19b)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9904[13:0] );

									end
									else
									if((r_sys_run_step==9'h19e)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9922[13:0] );

									end
									else
									if((r_sys_run_step==9'h199)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9892[13:0] );

									end
									else
									if((r_sys_run_step==9'h192)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9850[13:0] );

									end
									else
									if((r_sys_run_step==9'h197)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9880[13:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9802[13:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9820[13:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9826[13:0] );

									end
									else
									if((r_sys_run_step==9'h196)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9874[13:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9838[13:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9832[13:0] );

									end
									else
									if((r_sys_run_step==9'h198)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9886[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a0)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9934[13:0] );

									end
									else
									if((r_sys_run_step==9'h195)) begin
										r_sub18_T_addr <= $signed( w_sys_tmp9868[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h18b<=r_sys_run_step && r_sys_run_step<=9'h1a0)) begin
										r_sub18_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h18b<=r_sys_run_step && r_sys_run_step<=9'h1a0)) begin
										r_sub18_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h192)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5393[13:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5345[13:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5225[13:0] );

									end
									else
									if((r_sys_run_step==9'h188)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5273[13:0] );

									end
									else
									if((r_sys_run_step==9'h198)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5465[13:0] );

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5381[13:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5333[13:0] );

									end
									else
									if((r_sys_run_step==9'h196)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5441[13:0] );

									end
									else
									if((r_sys_run_step==9'h195)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5429[13:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5369[13:0] );

									end
									else
									if((r_sys_run_step==9'h199)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5477[13:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5321[13:0] );

									end
									else
									if((r_sys_run_step==9'h19a)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5489[13:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5357[13:0] );

									end
									else
									if((r_sys_run_step==9'h197)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5453[13:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5309[13:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5405[13:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5213[13:0] );

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5285[13:0] );

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5297[13:0] );

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5417[13:0] );

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_sub18_V_addr <= $signed( w_sys_tmp5261[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h185<=r_sys_run_step && r_sys_run_step<=9'h19a)) begin
										r_sub18_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h185<=r_sys_run_step && r_sys_run_step<=9'h19a)) begin
										r_sub18_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h192)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5393[13:0] );

									end
									else
									if((r_sys_run_step==9'h18e)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5345[13:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5225[13:0] );

									end
									else
									if((r_sys_run_step==9'h188)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5273[13:0] );

									end
									else
									if((r_sys_run_step==9'h198)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5465[13:0] );

									end
									else
									if((r_sys_run_step==9'h191)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5381[13:0] );

									end
									else
									if((r_sys_run_step==9'h18d)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5333[13:0] );

									end
									else
									if((r_sys_run_step==9'h196)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5441[13:0] );

									end
									else
									if((r_sys_run_step==9'h195)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5429[13:0] );

									end
									else
									if((r_sys_run_step==9'h190)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5369[13:0] );

									end
									else
									if((r_sys_run_step==9'h199)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5477[13:0] );

									end
									else
									if((r_sys_run_step==9'h18c)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5321[13:0] );

									end
									else
									if((r_sys_run_step==9'h19a)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5489[13:0] );

									end
									else
									if((r_sys_run_step==9'h18f)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5357[13:0] );

									end
									else
									if((r_sys_run_step==9'h197)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5453[13:0] );

									end
									else
									if((r_sys_run_step==9'h18b)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5309[13:0] );

									end
									else
									if((r_sys_run_step==9'h193)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5405[13:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5213[13:0] );

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5285[13:0] );

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5297[13:0] );

									end
									else
									if((r_sys_run_step==9'h194)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5417[13:0] );

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_sub18_U_addr <= $signed( w_sys_tmp5261[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h185<=r_sys_run_step && r_sys_run_step<=9'h19a)) begin
										r_sub18_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h185<=r_sys_run_step && r_sys_run_step<=9'h19a)) begin
										r_sub18_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12852[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12842[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12757[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12827[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12777[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12787[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12812[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12767[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12832[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12802[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12772[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12762[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12782[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12822[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12837[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12847[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12807[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12817[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12797[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub18_result_addr <= $signed( w_sys_tmp12792[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub18_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub18_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub18_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h4: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h63)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8032[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8020[13:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8086[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8038[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8068[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp7972[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8014[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp7990[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8002[13:0] );

									end
									else
									if((r_sys_run_step==9'h6b)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8080[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8074[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp7996[13:0] );

									end
									else
									if((r_sys_run_step==9'h6e)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8098[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8092[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8044[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8008[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8056[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8026[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp7966[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8050[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp8062[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h5a<=r_sys_run_step && r_sys_run_step<=9'h6e)) begin
										r_sub04_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h5a<=r_sys_run_step && r_sys_run_step<=9'h6e)) begin
										r_sub04_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6b)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1853[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1805[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1709[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1877[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1781[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1793[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1673[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1685[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1745[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1757[13:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1865[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1841[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1661[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1733[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1769[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1625[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1697[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1817[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1829[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1613[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp1721[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h59<=r_sys_run_step && r_sys_run_step<=9'h6d)) begin
										r_sub04_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h59<=r_sys_run_step && r_sys_run_step<=9'h6d)) begin
										r_sub04_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6b)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1853[13:0] );

									end
									else
									if((r_sys_run_step==9'h67)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1805[13:0] );

									end
									else
									if((r_sys_run_step==9'h5f)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1709[13:0] );

									end
									else
									if((r_sys_run_step==9'h6d)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1877[13:0] );

									end
									else
									if((r_sys_run_step==9'h65)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1781[13:0] );

									end
									else
									if((r_sys_run_step==9'h66)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1793[13:0] );

									end
									else
									if((r_sys_run_step==9'h5c)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1673[13:0] );

									end
									else
									if((r_sys_run_step==9'h5d)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1685[13:0] );

									end
									else
									if((r_sys_run_step==9'h62)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1745[13:0] );

									end
									else
									if((r_sys_run_step==9'h63)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1757[13:0] );

									end
									else
									if((r_sys_run_step==9'h6c)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1865[13:0] );

									end
									else
									if((r_sys_run_step==9'h6a)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1841[13:0] );

									end
									else
									if((r_sys_run_step==9'h5b)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1661[13:0] );

									end
									else
									if((r_sys_run_step==9'h61)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1733[13:0] );

									end
									else
									if((r_sys_run_step==9'h64)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1769[13:0] );

									end
									else
									if((r_sys_run_step==9'h5a)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1625[13:0] );

									end
									else
									if((r_sys_run_step==9'h5e)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1697[13:0] );

									end
									else
									if((r_sys_run_step==9'h68)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1817[13:0] );

									end
									else
									if((r_sys_run_step==9'h69)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1829[13:0] );

									end
									else
									if((r_sys_run_step==9'h59)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1613[13:0] );

									end
									else
									if((r_sys_run_step==9'h60)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp1721[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h59<=r_sys_run_step && r_sys_run_step<=9'h6d)) begin
										r_sub04_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h59<=r_sys_run_step && r_sys_run_step<=9'h6d)) begin
										r_sub04_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11447[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11417[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11382[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11412[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11452[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11392[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11407[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11437[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11377[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11422[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11402[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11362[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11457[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11387[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11432[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11427[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11397[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11372[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11462[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp11442[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h11: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub17_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub17_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h188)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9790[13:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9718[13:0] );

									end
									else
									if((r_sys_run_step==9'h182)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9754[13:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9670[13:0] );

									end
									else
									if((r_sys_run_step==9'h189)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9796[13:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9664[13:0] );

									end
									else
									if((r_sys_run_step==9'h181)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9748[13:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9724[13:0] );

									end
									else
									if((r_sys_run_step==9'h186)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9778[13:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9700[13:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9742[13:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9736[13:0] );

									end
									else
									if((r_sys_run_step==9'h18a)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9802[13:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9712[13:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9706[13:0] );

									end
									else
									if((r_sys_run_step==9'h185)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9772[13:0] );

									end
									else
									if((r_sys_run_step==9'h187)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9784[13:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9688[13:0] );

									end
									else
									if((r_sys_run_step==9'h184)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9766[13:0] );

									end
									else
									if((r_sys_run_step==9'h183)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9760[13:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9694[13:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_sub17_T_addr <= $signed( w_sys_tmp9730[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h175<=r_sys_run_step && r_sys_run_step<=9'h18a)) begin
										r_sub17_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h175<=r_sys_run_step && r_sys_run_step<=9'h18a)) begin
										r_sub17_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h171)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp4997[13:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp4949[13:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5105[13:0] );

									end
									else
									if((r_sys_run_step==9'h181)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5189[13:0] );

									end
									else
									if((r_sys_run_step==9'h184)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5225[13:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5069[13:0] );

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5033[13:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5081[13:0] );

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5021[13:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5141[13:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5045[13:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5129[13:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5117[13:0] );

									end
									else
									if((r_sys_run_step==9'h182)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5201[13:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5177[13:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5153[13:0] );

									end
									else
									if((r_sys_run_step==9'h183)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5213[13:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5165[13:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5057[13:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp4961[13:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5093[13:0] );

									end
									else
									if((r_sys_run_step==9'h172)) begin
										r_sub17_V_addr <= $signed( w_sys_tmp5009[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h16f<=r_sys_run_step && r_sys_run_step<=9'h184)) begin
										r_sub17_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h16f<=r_sys_run_step && r_sys_run_step<=9'h184)) begin
										r_sub17_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h171)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp4997[13:0] );

									end
									else
									if((r_sys_run_step==9'h16f)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp4949[13:0] );

									end
									else
									if((r_sys_run_step==9'h17a)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5105[13:0] );

									end
									else
									if((r_sys_run_step==9'h181)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5189[13:0] );

									end
									else
									if((r_sys_run_step==9'h184)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5225[13:0] );

									end
									else
									if((r_sys_run_step==9'h177)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5069[13:0] );

									end
									else
									if((r_sys_run_step==9'h174)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5033[13:0] );

									end
									else
									if((r_sys_run_step==9'h178)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5081[13:0] );

									end
									else
									if((r_sys_run_step==9'h173)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5021[13:0] );

									end
									else
									if((r_sys_run_step==9'h17d)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5141[13:0] );

									end
									else
									if((r_sys_run_step==9'h175)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5045[13:0] );

									end
									else
									if((r_sys_run_step==9'h17c)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5129[13:0] );

									end
									else
									if((r_sys_run_step==9'h17b)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5117[13:0] );

									end
									else
									if((r_sys_run_step==9'h182)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5201[13:0] );

									end
									else
									if((r_sys_run_step==9'h180)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5177[13:0] );

									end
									else
									if((r_sys_run_step==9'h17e)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5153[13:0] );

									end
									else
									if((r_sys_run_step==9'h183)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5213[13:0] );

									end
									else
									if((r_sys_run_step==9'h17f)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5165[13:0] );

									end
									else
									if((r_sys_run_step==9'h176)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5057[13:0] );

									end
									else
									if((r_sys_run_step==9'h170)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp4961[13:0] );

									end
									else
									if((r_sys_run_step==9'h179)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5093[13:0] );

									end
									else
									if((r_sys_run_step==9'h172)) begin
										r_sub17_U_addr <= $signed( w_sys_tmp5009[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h16f<=r_sys_run_step && r_sys_run_step<=9'h184)) begin
										r_sub17_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h16f<=r_sys_run_step && r_sys_run_step<=9'h184)) begin
										r_sub17_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12697[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12742[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12677[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12722[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12737[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12702[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12747[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12682[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12727[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12707[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12662[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12687[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12712[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12667[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12732[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12672[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12717[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12752[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12692[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_addr <= $signed( w_sys_tmp12657[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub17_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub17_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub17_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'ha: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub10_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub10_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he8)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8830[13:0] );

									end
									else
									if((r_sys_run_step==9'hf0)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8878[13:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8824[13:0] );

									end
									else
									if((r_sys_run_step==9'hef)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8872[13:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8818[13:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8794[13:0] );

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8854[13:0] );

									end
									else
									if((r_sys_run_step==9'hf1)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8884[13:0] );

									end
									else
									if((r_sys_run_step==9'hee)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8866[13:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8758[13:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8782[13:0] );

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8842[13:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8836[13:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8776[13:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8806[13:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8800[13:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8770[13:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8812[13:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8788[13:0] );

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8860[13:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8764[13:0] );

									end
									else
									if((r_sys_run_step==9'heb)) begin
										r_sub10_T_addr <= $signed( w_sys_tmp8848[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hdc<=r_sys_run_step && r_sys_run_step<=9'hf1)) begin
										r_sub10_T_datain <= w_sys_tmp7452;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hdc<=r_sys_run_step && r_sys_run_step<=9'hf1)) begin
										r_sub10_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd9)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3173[13:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3329[13:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3305[13:0] );

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3413[13:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3353[13:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3341[13:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3197[13:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3293[13:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3281[13:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3365[13:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3245[13:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3317[13:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3221[13:0] );

									end
									else
									if((r_sys_run_step==9'heb)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3389[13:0] );

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3401[13:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3209[13:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3257[13:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3185[13:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3233[13:0] );

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3377[13:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_sub10_V_addr <= $signed( w_sys_tmp3269[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hd9<=r_sys_run_step && r_sys_run_step<=9'hed)) begin
										r_sub10_V_datain <= w_sys_tmp601;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hd9<=r_sys_run_step && r_sys_run_step<=9'hed)) begin
										r_sub10_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd9)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3173[13:0] );

									end
									else
									if((r_sys_run_step==9'he6)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3329[13:0] );

									end
									else
									if((r_sys_run_step==9'he4)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3305[13:0] );

									end
									else
									if((r_sys_run_step==9'hed)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3413[13:0] );

									end
									else
									if((r_sys_run_step==9'he8)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3353[13:0] );

									end
									else
									if((r_sys_run_step==9'he7)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3341[13:0] );

									end
									else
									if((r_sys_run_step==9'hdb)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3197[13:0] );

									end
									else
									if((r_sys_run_step==9'he3)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3293[13:0] );

									end
									else
									if((r_sys_run_step==9'he2)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3281[13:0] );

									end
									else
									if((r_sys_run_step==9'he9)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3365[13:0] );

									end
									else
									if((r_sys_run_step==9'hdf)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3245[13:0] );

									end
									else
									if((r_sys_run_step==9'he5)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3317[13:0] );

									end
									else
									if((r_sys_run_step==9'hdd)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3221[13:0] );

									end
									else
									if((r_sys_run_step==9'heb)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3389[13:0] );

									end
									else
									if((r_sys_run_step==9'hec)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3401[13:0] );

									end
									else
									if((r_sys_run_step==9'hdc)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3209[13:0] );

									end
									else
									if((r_sys_run_step==9'he0)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3257[13:0] );

									end
									else
									if((r_sys_run_step==9'hda)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3185[13:0] );

									end
									else
									if((r_sys_run_step==9'hde)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3233[13:0] );

									end
									else
									if((r_sys_run_step==9'hea)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3377[13:0] );

									end
									else
									if((r_sys_run_step==9'he1)) begin
										r_sub10_U_addr <= $signed( w_sys_tmp3269[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hd9<=r_sys_run_step && r_sys_run_step<=9'hed)) begin
										r_sub10_U_datain <= w_sys_tmp595;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'hd9<=r_sys_run_step && r_sys_run_step<=9'hed)) begin
										r_sub10_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp11962[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp11987[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12052[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp11977[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12007[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp11982[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12022[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12027[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12047[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp11972[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12037[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp11967[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12057[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12042[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp11997[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12017[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12032[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp11992[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12002[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub10_result_addr <= $signed( w_sys_tmp12012[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub10_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub10_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub10_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h14: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub20_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub20_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10198[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10096[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10168[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10144[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10120[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10192[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10150[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10078[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10126[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10084[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10162[13:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10186[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10132[13:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10180[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10174[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10102[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10072[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10090[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10114[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10156[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10138[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub20_T_addr <= $signed( w_sys_tmp10108[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h17)) begin
										r_sub20_T_datain <= w_sys_tmp10074;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h17)) begin
										r_sub20_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5783[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5891[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5771[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5843[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5903[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5951[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5939[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5807[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5759[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5855[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5867[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5831[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5795[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5879[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5915[13:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5975[13:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5987[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5963[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5927[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5819[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub20_V_addr <= $signed( w_sys_tmp5999[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h16)) begin
										r_sub20_V_datain <= w_sys_tmp5767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h16)) begin
										r_sub20_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5783[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5891[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5771[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5843[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5903[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5951[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5939[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5807[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5759[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5855[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5867[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5831[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5795[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5879[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5915[13:0] );

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5975[13:0] );

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5987[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5963[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5927[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5819[13:0] );

									end
									else
									if((r_sys_run_step==9'h16)) begin
										r_sub20_U_addr <= $signed( w_sys_tmp5999[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h16)) begin
										r_sub20_U_datain <= w_sys_tmp5761;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h2<=r_sys_run_step && r_sys_run_step<=9'h16)) begin
										r_sub20_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13060[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13030[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp12964[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13018[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13042[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13000[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13048[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13066[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13054[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp12988[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13006[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp12976[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp12982[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp12994[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13036[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp12970[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13024[13:0] );

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13072[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp12958[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub20_result_addr <= $signed( w_sys_tmp13012[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub20_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub20_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub20_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h15: begin
									if((r_sys_run_step==9'h1)) begin
										r_sub21_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub21_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10198[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10228[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10318[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10240[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10258[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10192[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10312[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10222[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10300[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10264[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10270[13:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10324[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10288[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10306[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10276[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10246[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10216[13:0] );

									end
									else
									if((r_sys_run_step==9'h27)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10294[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10252[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10282[13:0] );

									end
									else
									if((r_sys_run_step==9'h2d)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10330[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub21_T_addr <= $signed( w_sys_tmp10234[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h18<=r_sys_run_step && r_sys_run_step<=9'h2d)) begin
										r_sub21_T_datain <= w_sys_tmp10074;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h18<=r_sys_run_step && r_sys_run_step<=9'h2d)) begin
										r_sub21_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_V_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h27)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6203[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6107[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6155[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6095[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6047[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6167[13:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6263[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6191[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6059[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6239[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6215[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6083[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6179[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6071[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6251[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6035[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6023[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6131[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6143[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6227[13:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp5999[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub21_V_addr <= $signed( w_sys_tmp6119[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h17<=r_sys_run_step && r_sys_run_step<=9'h2c)) begin
										r_sub21_V_datain <= w_sys_tmp5767;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h17<=r_sys_run_step && r_sys_run_step<=9'h2c)) begin
										r_sub21_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h27)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6203[13:0] );

									end
									else
									if((r_sys_run_step==9'h1f)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6107[13:0] );

									end
									else
									if((r_sys_run_step==9'h23)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6155[13:0] );

									end
									else
									if((r_sys_run_step==9'h1e)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6095[13:0] );

									end
									else
									if((r_sys_run_step==9'h1a)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6047[13:0] );

									end
									else
									if((r_sys_run_step==9'h24)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6167[13:0] );

									end
									else
									if((r_sys_run_step==9'h2c)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6263[13:0] );

									end
									else
									if((r_sys_run_step==9'h26)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6191[13:0] );

									end
									else
									if((r_sys_run_step==9'h1b)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6059[13:0] );

									end
									else
									if((r_sys_run_step==9'h2a)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6239[13:0] );

									end
									else
									if((r_sys_run_step==9'h28)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6215[13:0] );

									end
									else
									if((r_sys_run_step==9'h1d)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6083[13:0] );

									end
									else
									if((r_sys_run_step==9'h25)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6179[13:0] );

									end
									else
									if((r_sys_run_step==9'h1c)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6071[13:0] );

									end
									else
									if((r_sys_run_step==9'h2b)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6251[13:0] );

									end
									else
									if((r_sys_run_step==9'h19)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6035[13:0] );

									end
									else
									if((r_sys_run_step==9'h18)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6023[13:0] );

									end
									else
									if((r_sys_run_step==9'h21)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6131[13:0] );

									end
									else
									if((r_sys_run_step==9'h22)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6143[13:0] );

									end
									else
									if((r_sys_run_step==9'h29)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6227[13:0] );

									end
									else
									if((r_sys_run_step==9'h17)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp5999[13:0] );

									end
									else
									if((r_sys_run_step==9'h20)) begin
										r_sub21_U_addr <= $signed( w_sys_tmp6119[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h17<=r_sys_run_step && r_sys_run_step<=9'h2c)) begin
										r_sub21_U_datain <= w_sys_tmp5761;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h17<=r_sys_run_step && r_sys_run_step<=9'h2c)) begin
										r_sub21_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_addr <= 14'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13173[13:0] );

									end
									else
									if((r_sys_run_step==9'h8)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13118[13:0] );

									end
									else
									if((r_sys_run_step==9'h9)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13123[13:0] );

									end
									else
									if((r_sys_run_step==9'he)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13148[13:0] );

									end
									else
									if((r_sys_run_step==9'h1)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13083[13:0] );

									end
									else
									if((r_sys_run_step==9'h6)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13108[13:0] );

									end
									else
									if((r_sys_run_step==9'ha)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13128[13:0] );

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13163[13:0] );

									end
									else
									if((r_sys_run_step==9'h7)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13113[13:0] );

									end
									else
									if((r_sys_run_step==9'hb)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13133[13:0] );

									end
									else
									if((r_sys_run_step==9'h5)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13103[13:0] );

									end
									else
									if((r_sys_run_step==9'hd)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13143[13:0] );

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13158[13:0] );

									end
									else
									if((r_sys_run_step==9'h3)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13093[13:0] );

									end
									else
									if((r_sys_run_step==9'hc)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13138[13:0] );

									end
									else
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13078[13:0] );

									end
									else
									if((r_sys_run_step==9'hf)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13153[13:0] );

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13168[13:0] );

									end
									else
									if((r_sys_run_step==9'h2)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13088[13:0] );

									end
									else
									if((r_sys_run_step==9'h4)) begin
										r_sub21_result_addr <= $signed( w_sys_tmp13098[13:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub21_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h1: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h2: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h3: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h4: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h5: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h6: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h7: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h8: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h9: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'ha: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hb: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hc: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hd: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'he: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'hf: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h10: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h11: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h12: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h13: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h14: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h15: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h16: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h17: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

								5'h18: begin
									if((r_sys_run_step==9'h0)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((9'h0<=r_sys_run_step && r_sys_run_step<=9'h13)) begin
										r_sub21_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub21_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp0_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h23)) begin
										r_sys_tmp0_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp1_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h22)) begin
										r_sys_tmp1_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp2_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h21)) begin
										r_sys_tmp2_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp3_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h20)) begin
										r_sys_tmp3_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1f)) begin
										r_sys_tmp4_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11) || (r_sys_run_step==9'h17)) begin
										r_sys_tmp5_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1e)) begin
										r_sys_tmp5_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h2f)) begin
										r_sys_tmp6_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1d)) begin
										r_sys_tmp6_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he) || (r_sys_run_step==9'h10) || (r_sys_run_step==9'h14)) begin
										r_sys_tmp7_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1c)) begin
										r_sys_tmp7_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19) || (r_sys_run_step==9'h21) || (r_sys_run_step==9'h2a) || (r_sys_run_step==9'h33)) begin
										r_sys_tmp8_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1b)) begin
										r_sys_tmp8_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17) || (r_sys_run_step==9'h1e) || (r_sys_run_step==9'h27) || (r_sys_run_step==9'h30)) begin
										r_sys_tmp9_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h1a)) begin
										r_sys_tmp9_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14) || (r_sys_run_step==9'h18) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h32)) begin
										r_sys_tmp10_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h19)) begin
										r_sys_tmp10_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h29) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h3c)) begin
										r_sys_tmp11_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h18)) begin
										r_sys_tmp11_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc) || (r_sys_run_step==9'hd) || (r_sys_run_step==9'hf) || (r_sys_run_step==9'h12) || (r_sys_run_step==9'h19)) begin
										r_sys_tmp12_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h17)) begin
										r_sys_tmp12_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h32) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h40)) begin
										r_sys_tmp13_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp13_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12) || (r_sys_run_step==9'h15) || (r_sys_run_step==9'h1c) || (r_sys_run_step==9'h24) || (r_sys_run_step==9'h2d) || (r_sys_run_step==9'h38)) begin
										r_sys_tmp14_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h16)) begin
										r_sys_tmp14_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h20) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h38) || (r_sys_run_step==9'h3e)) begin
										r_sys_tmp15_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp15_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10) || (r_sys_run_step==9'h13) || (r_sys_run_step==9'h1a) || (r_sys_run_step==9'h23) || (r_sys_run_step==9'h2c) || (r_sys_run_step==9'h35) || (r_sys_run_step==9'h3a) || (r_sys_run_step==9'h3e)) begin
										r_sys_tmp16_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp16_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf) || (r_sys_run_step==9'h11) || (r_sys_run_step==9'h16) || (r_sys_run_step==9'h1d) || (r_sys_run_step==9'h26) || (r_sys_run_step==9'h2f) || (r_sys_run_step==9'h36) || (r_sys_run_step==9'h3c) || (r_sys_run_step==9'h40)) begin
										r_sys_tmp17_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp17_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp18_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp18_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp19_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp19_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp20_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp20_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp21_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp21_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp22_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp22_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp23_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp23_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp24_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp24_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp25_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp25_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp26_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp26_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp27_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp27_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp28_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp28_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp29_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp29_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp30_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp30_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp31_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp31_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp32_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp32_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp33_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp33_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp34_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp34_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp35_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp35_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp36_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp36_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp37_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp37_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp38_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp38_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp39_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp39_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp40_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp40_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp41_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp41_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp42_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp42_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp43_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp43_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp44_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp44_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp45_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp45_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp46_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp46_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp47_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp47_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp48_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp48_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp49_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp49_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp50_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp50_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp51_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp51_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp52_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp52_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp53_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp53_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp54_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp54_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp55_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp55_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp56_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp56_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp57_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp57_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp58_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp58_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp59_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp59_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp60_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp60_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp61_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp61_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp62_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp62_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp63_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp63_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp64_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp64_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp65_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp65_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp66_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp66_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp67_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp67_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp68_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp68_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp69_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp69_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp70_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp70_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp71_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp71_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp72_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp72_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp73_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp73_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp74_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp74_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp75_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp75_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp76_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp76_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp77_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp77_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp78_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp78_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp79_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp79_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp80_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp80_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp81_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp81_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp82_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp82_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp83_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp83_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp84_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp84_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp85_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp85_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp86_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp86_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp87_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp87_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp88_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp88_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp89_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp89_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp90_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp90_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp91_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp91_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp92_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp92_float <= w_sub21_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp93_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp93_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp94_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp94_float <= w_sub23_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp95_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp95_float <= w_sub24_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp96_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp97_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp98_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp99_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp100_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp101_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp102_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp102_float <= w_sub22_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp103_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp104_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp105_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp106_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp107_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp108_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp109_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp110_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp111_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp112_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp113_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp114_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp115_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp116_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp117_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp118_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp119_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp120_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp121_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp122_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp123_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp124_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp125_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp126_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp127_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp128_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp129_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp130_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp131_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp132_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp133_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp134_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp135_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp136_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf)) begin
										r_sys_tmp137_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp138_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp139_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp140_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp141_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp142_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp143_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp144_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp145_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp146_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp147_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp148_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp149_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp150_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp151_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp152_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp153_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp154_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he)) begin
										r_sys_tmp155_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp156_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp157_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp158_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp159_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp160_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp161_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp162_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp163_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp164_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp165_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp166_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp167_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp168_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp169_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp170_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp171_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp172_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd)) begin
										r_sys_tmp173_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp174_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp175_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp176_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp177_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp178_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp179_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp180_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp181_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp182_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp183_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp184_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp185_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp186_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp187_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp188_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp189_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp190_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc)) begin
										r_sys_tmp191_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp192_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp193_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp194_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp195_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp196_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp197_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp198_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp199_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp200_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp201_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp202_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp203_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp204_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp205_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp206_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp207_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp208_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb)) begin
										r_sys_tmp209_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp210_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp211_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp212_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp213_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp214_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp215_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp216_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp217_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp218_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp219_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp220_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp221_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp222_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp223_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp224_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp225_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp226_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha)) begin
										r_sys_tmp227_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp228_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp229_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp230_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp231_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp232_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp233_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp234_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp235_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp236_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp237_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp238_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp239_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp240_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp241_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp242_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp243_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp244_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h9)) begin
										r_sys_tmp245_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp246_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp247_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp248_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp249_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp250_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp251_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp252_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp253_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp254_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp255_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp256_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp257_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp258_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp259_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp260_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp261_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp262_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h8)) begin
										r_sys_tmp263_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp264_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp265_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp266_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp267_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp268_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp269_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp270_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp271_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp272_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp273_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp274_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp275_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp276_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp277_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp278_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp279_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp280_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h7)) begin
										r_sys_tmp281_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp282_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp283_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp284_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp285_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp286_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp287_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp288_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp289_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp290_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp291_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp292_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp293_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp294_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp295_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp296_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp297_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp298_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h6)) begin
										r_sys_tmp299_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp300_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp301_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp302_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp303_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp304_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp305_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp306_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp307_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp308_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp309_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp310_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp311_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp312_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp313_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp314_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp315_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp316_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h5)) begin
										r_sys_tmp317_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp318_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp319_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp320_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp321_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp322_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp323_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp324_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp325_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp326_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp327_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp328_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp329_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp330_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp331_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp332_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp333_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp334_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h4)) begin
										r_sys_tmp335_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp336_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp337_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp338_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp339_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp340_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp341_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp342_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp343_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp344_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp345_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp346_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp347_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp348_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp349_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp350_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp351_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp352_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h3)) begin
										r_sys_tmp353_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp354_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp355_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp356_float <= w_sub09_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp357_float <= w_sub12_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp358_float <= w_sub15_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp359_float <= w_sub17_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp360_float <= w_sub19_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp361_float <= w_sub18_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp362_float <= w_sub16_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp363_float <= w_sub14_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp364_float <= w_sub13_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp365_float <= w_sub11_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp366_float <= w_sub10_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp367_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp368_float <= w_sub06_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp369_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp370_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2)) begin
										r_sys_tmp371_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hf) || (r_sys_run_step==9'h23)) begin
										r_sys_tmp372_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'he) || (r_sys_run_step==9'h22)) begin
										r_sys_tmp373_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hd) || (r_sys_run_step==9'h21)) begin
										r_sys_tmp374_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hc) || (r_sys_run_step==9'h20)) begin
										r_sys_tmp375_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'hb) || (r_sys_run_step==9'h1f)) begin
										r_sys_tmp376_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'ha) || (r_sys_run_step==9'h1e)) begin
										r_sys_tmp377_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h29)) begin
										r_sys_tmp378_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h15)) begin
										r_sys_tmp378_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h28)) begin
										r_sys_tmp379_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h14)) begin
										r_sys_tmp379_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h27)) begin
										r_sys_tmp380_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h13)) begin
										r_sys_tmp380_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h26)) begin
										r_sys_tmp381_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h12)) begin
										r_sys_tmp381_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h25)) begin
										r_sys_tmp382_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h11)) begin
										r_sys_tmp382_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h24)) begin
										r_sys_tmp383_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h10)) begin
										r_sys_tmp383_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h31)) begin
										r_sys_tmp384_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h9) || (r_sys_run_step==9'h1d)) begin
										r_sys_tmp384_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h30)) begin
										r_sys_tmp385_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h8) || (r_sys_run_step==9'h1c)) begin
										r_sys_tmp385_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2f)) begin
										r_sys_tmp386_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h7) || (r_sys_run_step==9'h1b)) begin
										r_sys_tmp386_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2e)) begin
										r_sys_tmp387_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h6) || (r_sys_run_step==9'h1a)) begin
										r_sys_tmp387_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2d)) begin
										r_sys_tmp388_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h5) || (r_sys_run_step==9'h19)) begin
										r_sys_tmp388_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2c)) begin
										r_sys_tmp389_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h4) || (r_sys_run_step==9'h18)) begin
										r_sys_tmp389_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2b)) begin
										r_sys_tmp390_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h3) || (r_sys_run_step==9'h17)) begin
										r_sys_tmp390_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								5'h0: begin
									if((r_sys_run_step==9'h2a)) begin
										r_sys_tmp391_float <= w_sub02_result_dataout;

									end
									else
									if((r_sys_run_step==9'h2) || (r_sys_run_step==9'h16)) begin
										r_sys_tmp391_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
