/*
TimeStamp:	2016/6/26		17:47
*/


module P3_2dim(
	input                 clock,	
	input                 reset_n,	
	input                 ce,	
	input                 i_run_req,	
	output                o_run_busy	
);

	reg         [31:0] r_ip_AddFloat_portA_0;
	reg         [31:0] r_ip_AddFloat_portB_0;
	wire        [31:0] w_ip_AddFloat_result_0;
	reg         [31:0] r_ip_MultFloat_multiplicand_0;
	reg         [31:0] r_ip_MultFloat_multiplier_0;
	wire        [31:0] w_ip_MultFloat_product_0;
	reg  signed [31:0] r_ip_FixedToFloat_fixed_0;
	wire        [31:0] w_ip_FixedToFloat_floating_0;
	reg         [ 1:0] r_sys_processing_methodID;
	wire               w_sys_boolTrue;
	wire               w_sys_boolFalse;
	wire signed [31:0] w_sys_intOne;
	wire signed [31:0] w_sys_intZero;
	wire               w_sys_ce;
	reg         [ 1:0] r_sys_run_caller;
	reg                r_sys_run_req;
	reg         [ 6:0] r_sys_run_phase;
	reg         [ 3:0] r_sys_run_stage;
	reg         [ 6:0] r_sys_run_step;
	reg                r_sys_run_busy;
	wire        [ 3:0] w_sys_run_stage_p1;
	wire        [ 6:0] w_sys_run_step_p1;
	wire signed [ 8:0] w_fld_T_0_addr_0;
	wire        [31:0] w_fld_T_0_datain_0;
	wire        [31:0] w_fld_T_0_dataout_0;
	wire               w_fld_T_0_r_w_0;
	wire               w_fld_T_0_ce_0;
	reg  signed [ 8:0] r_fld_T_0_addr_1;
	reg         [31:0] r_fld_T_0_datain_1;
	wire        [31:0] w_fld_T_0_dataout_1;
	reg                r_fld_T_0_r_w_1;
	wire               w_fld_T_0_ce_1;
	wire signed [ 8:0] w_fld_TT_1_addr_0;
	wire        [31:0] w_fld_TT_1_datain_0;
	wire        [31:0] w_fld_TT_1_dataout_0;
	wire               w_fld_TT_1_r_w_0;
	wire               w_fld_TT_1_ce_0;
	reg  signed [ 8:0] r_fld_TT_1_addr_1;
	reg         [31:0] r_fld_TT_1_datain_1;
	wire        [31:0] w_fld_TT_1_dataout_1;
	reg                r_fld_TT_1_r_w_1;
	wire               w_fld_TT_1_ce_1;
	wire signed [ 8:0] w_fld_U_2_addr_0;
	wire        [31:0] w_fld_U_2_datain_0;
	wire        [31:0] w_fld_U_2_dataout_0;
	wire               w_fld_U_2_r_w_0;
	wire               w_fld_U_2_ce_0;
	reg  signed [ 8:0] r_fld_U_2_addr_1;
	reg         [31:0] r_fld_U_2_datain_1;
	wire        [31:0] w_fld_U_2_dataout_1;
	reg                r_fld_U_2_r_w_1;
	wire               w_fld_U_2_ce_1;
	wire signed [ 8:0] w_fld_V_3_addr_0;
	wire        [31:0] w_fld_V_3_datain_0;
	wire        [31:0] w_fld_V_3_dataout_0;
	wire               w_fld_V_3_r_w_0;
	wire               w_fld_V_3_ce_0;
	reg  signed [ 8:0] r_fld_V_3_addr_1;
	reg         [31:0] r_fld_V_3_datain_1;
	wire        [31:0] w_fld_V_3_dataout_1;
	reg                r_fld_V_3_r_w_1;
	wire               w_fld_V_3_ce_1;
	reg  signed [31:0] r_run_k_13;
	reg  signed [31:0] r_run_j_14;
	reg  signed [31:0] r_run_n_15;
	reg  signed [31:0] r_run_mx_16;
	reg  signed [31:0] r_run_my_17;
	reg         [31:0] r_run_dt_18;
	reg         [31:0] r_run_dx_19;
	reg         [31:0] r_run_dy_20;
	reg         [31:0] r_run_r1_21;
	reg         [31:0] r_run_r2_22;
	reg         [31:0] r_run_r3_23;
	reg         [31:0] r_run_r4_24;
	reg         [31:0] r_run_YY_25;
	reg  signed [31:0] r_run_kx_26;
	reg  signed [31:0] r_run_ky_27;
	reg  signed [31:0] r_run_nlast_28;
	reg  signed [31:0] r_run_copy0_j_29;
	reg  signed [31:0] r_run_copy1_j_30;
	reg  signed [31:0] r_run_copy2_j_31;
	reg  signed [31:0] r_run_copy0_j_32;
	reg                r_sub08_run_req;
	wire               w_sub08_run_busy;
	wire signed [ 9:0] w_sub08_T_addr;
	reg  signed [ 9:0] r_sub08_T_addr;
	wire        [31:0] w_sub08_T_datain;
	reg         [31:0] r_sub08_T_datain;
	wire        [31:0] w_sub08_T_dataout;
	wire               w_sub08_T_r_w;
	reg                r_sub08_T_r_w;
	wire signed [ 9:0] w_sub08_V_addr;
	reg  signed [ 9:0] r_sub08_V_addr;
	wire        [31:0] w_sub08_V_datain;
	reg         [31:0] r_sub08_V_datain;
	wire        [31:0] w_sub08_V_dataout;
	wire               w_sub08_V_r_w;
	reg                r_sub08_V_r_w;
	wire signed [ 9:0] w_sub08_U_addr;
	reg  signed [ 9:0] r_sub08_U_addr;
	wire        [31:0] w_sub08_U_datain;
	reg         [31:0] r_sub08_U_datain;
	wire        [31:0] w_sub08_U_dataout;
	wire               w_sub08_U_r_w;
	reg                r_sub08_U_r_w;
	wire signed [ 9:0] w_sub08_result_addr;
	reg  signed [ 9:0] r_sub08_result_addr;
	wire        [31:0] w_sub08_result_datain;
	reg         [31:0] r_sub08_result_datain;
	wire        [31:0] w_sub08_result_dataout;
	wire               w_sub08_result_r_w;
	reg                r_sub08_result_r_w;
	reg                r_sub03_run_req;
	wire               w_sub03_run_busy;
	wire signed [ 9:0] w_sub03_T_addr;
	reg  signed [ 9:0] r_sub03_T_addr;
	wire        [31:0] w_sub03_T_datain;
	reg         [31:0] r_sub03_T_datain;
	wire        [31:0] w_sub03_T_dataout;
	wire               w_sub03_T_r_w;
	reg                r_sub03_T_r_w;
	wire signed [ 9:0] w_sub03_V_addr;
	reg  signed [ 9:0] r_sub03_V_addr;
	wire        [31:0] w_sub03_V_datain;
	reg         [31:0] r_sub03_V_datain;
	wire        [31:0] w_sub03_V_dataout;
	wire               w_sub03_V_r_w;
	reg                r_sub03_V_r_w;
	wire signed [ 9:0] w_sub03_U_addr;
	reg  signed [ 9:0] r_sub03_U_addr;
	wire        [31:0] w_sub03_U_datain;
	reg         [31:0] r_sub03_U_datain;
	wire        [31:0] w_sub03_U_dataout;
	wire               w_sub03_U_r_w;
	reg                r_sub03_U_r_w;
	wire signed [ 9:0] w_sub03_result_addr;
	reg  signed [ 9:0] r_sub03_result_addr;
	wire        [31:0] w_sub03_result_datain;
	reg         [31:0] r_sub03_result_datain;
	wire        [31:0] w_sub03_result_dataout;
	wire               w_sub03_result_r_w;
	reg                r_sub03_result_r_w;
	reg                r_sub02_run_req;
	wire               w_sub02_run_busy;
	wire signed [ 9:0] w_sub02_T_addr;
	reg  signed [ 9:0] r_sub02_T_addr;
	wire        [31:0] w_sub02_T_datain;
	reg         [31:0] r_sub02_T_datain;
	wire        [31:0] w_sub02_T_dataout;
	wire               w_sub02_T_r_w;
	reg                r_sub02_T_r_w;
	wire signed [ 9:0] w_sub02_V_addr;
	reg  signed [ 9:0] r_sub02_V_addr;
	wire        [31:0] w_sub02_V_datain;
	reg         [31:0] r_sub02_V_datain;
	wire        [31:0] w_sub02_V_dataout;
	wire               w_sub02_V_r_w;
	reg                r_sub02_V_r_w;
	wire signed [ 9:0] w_sub02_U_addr;
	reg  signed [ 9:0] r_sub02_U_addr;
	wire        [31:0] w_sub02_U_datain;
	reg         [31:0] r_sub02_U_datain;
	wire        [31:0] w_sub02_U_dataout;
	wire               w_sub02_U_r_w;
	reg                r_sub02_U_r_w;
	wire signed [ 9:0] w_sub02_result_addr;
	reg  signed [ 9:0] r_sub02_result_addr;
	wire        [31:0] w_sub02_result_datain;
	reg         [31:0] r_sub02_result_datain;
	wire        [31:0] w_sub02_result_dataout;
	wire               w_sub02_result_r_w;
	reg                r_sub02_result_r_w;
	reg                r_sub01_run_req;
	wire               w_sub01_run_busy;
	wire signed [ 9:0] w_sub01_T_addr;
	reg  signed [ 9:0] r_sub01_T_addr;
	wire        [31:0] w_sub01_T_datain;
	reg         [31:0] r_sub01_T_datain;
	wire        [31:0] w_sub01_T_dataout;
	wire               w_sub01_T_r_w;
	reg                r_sub01_T_r_w;
	wire signed [ 9:0] w_sub01_V_addr;
	reg  signed [ 9:0] r_sub01_V_addr;
	wire        [31:0] w_sub01_V_datain;
	reg         [31:0] r_sub01_V_datain;
	wire        [31:0] w_sub01_V_dataout;
	wire               w_sub01_V_r_w;
	reg                r_sub01_V_r_w;
	wire signed [ 9:0] w_sub01_U_addr;
	reg  signed [ 9:0] r_sub01_U_addr;
	wire        [31:0] w_sub01_U_datain;
	reg         [31:0] r_sub01_U_datain;
	wire        [31:0] w_sub01_U_dataout;
	wire               w_sub01_U_r_w;
	reg                r_sub01_U_r_w;
	wire signed [ 9:0] w_sub01_result_addr;
	reg  signed [ 9:0] r_sub01_result_addr;
	wire        [31:0] w_sub01_result_datain;
	reg         [31:0] r_sub01_result_datain;
	wire        [31:0] w_sub01_result_dataout;
	wire               w_sub01_result_r_w;
	reg                r_sub01_result_r_w;
	reg                r_sub00_run_req;
	wire               w_sub00_run_busy;
	wire signed [ 9:0] w_sub00_T_addr;
	reg  signed [ 9:0] r_sub00_T_addr;
	wire        [31:0] w_sub00_T_datain;
	reg         [31:0] r_sub00_T_datain;
	wire        [31:0] w_sub00_T_dataout;
	wire               w_sub00_T_r_w;
	reg                r_sub00_T_r_w;
	wire signed [ 9:0] w_sub00_V_addr;
	reg  signed [ 9:0] r_sub00_V_addr;
	wire        [31:0] w_sub00_V_datain;
	reg         [31:0] r_sub00_V_datain;
	wire        [31:0] w_sub00_V_dataout;
	wire               w_sub00_V_r_w;
	reg                r_sub00_V_r_w;
	wire signed [ 9:0] w_sub00_U_addr;
	reg  signed [ 9:0] r_sub00_U_addr;
	wire        [31:0] w_sub00_U_datain;
	reg         [31:0] r_sub00_U_datain;
	wire        [31:0] w_sub00_U_dataout;
	wire               w_sub00_U_r_w;
	reg                r_sub00_U_r_w;
	wire signed [ 9:0] w_sub00_result_addr;
	reg  signed [ 9:0] r_sub00_result_addr;
	wire        [31:0] w_sub00_result_datain;
	reg         [31:0] r_sub00_result_datain;
	wire        [31:0] w_sub00_result_dataout;
	wire               w_sub00_result_r_w;
	reg                r_sub00_result_r_w;
	reg                r_sub07_run_req;
	wire               w_sub07_run_busy;
	wire signed [ 9:0] w_sub07_T_addr;
	reg  signed [ 9:0] r_sub07_T_addr;
	wire        [31:0] w_sub07_T_datain;
	reg         [31:0] r_sub07_T_datain;
	wire        [31:0] w_sub07_T_dataout;
	wire               w_sub07_T_r_w;
	reg                r_sub07_T_r_w;
	wire signed [ 9:0] w_sub07_V_addr;
	reg  signed [ 9:0] r_sub07_V_addr;
	wire        [31:0] w_sub07_V_datain;
	reg         [31:0] r_sub07_V_datain;
	wire        [31:0] w_sub07_V_dataout;
	wire               w_sub07_V_r_w;
	reg                r_sub07_V_r_w;
	wire signed [ 9:0] w_sub07_U_addr;
	reg  signed [ 9:0] r_sub07_U_addr;
	wire        [31:0] w_sub07_U_datain;
	reg         [31:0] r_sub07_U_datain;
	wire        [31:0] w_sub07_U_dataout;
	wire               w_sub07_U_r_w;
	reg                r_sub07_U_r_w;
	wire signed [ 9:0] w_sub07_result_addr;
	reg  signed [ 9:0] r_sub07_result_addr;
	wire        [31:0] w_sub07_result_datain;
	reg         [31:0] r_sub07_result_datain;
	wire        [31:0] w_sub07_result_dataout;
	wire               w_sub07_result_r_w;
	reg                r_sub07_result_r_w;
	reg                r_sub06_run_req;
	wire               w_sub06_run_busy;
	wire signed [ 9:0] w_sub06_T_addr;
	reg  signed [ 9:0] r_sub06_T_addr;
	wire        [31:0] w_sub06_T_datain;
	reg         [31:0] r_sub06_T_datain;
	wire        [31:0] w_sub06_T_dataout;
	wire               w_sub06_T_r_w;
	reg                r_sub06_T_r_w;
	wire signed [ 9:0] w_sub06_V_addr;
	reg  signed [ 9:0] r_sub06_V_addr;
	wire        [31:0] w_sub06_V_datain;
	reg         [31:0] r_sub06_V_datain;
	wire        [31:0] w_sub06_V_dataout;
	wire               w_sub06_V_r_w;
	reg                r_sub06_V_r_w;
	wire signed [ 9:0] w_sub06_U_addr;
	reg  signed [ 9:0] r_sub06_U_addr;
	wire        [31:0] w_sub06_U_datain;
	reg         [31:0] r_sub06_U_datain;
	wire        [31:0] w_sub06_U_dataout;
	wire               w_sub06_U_r_w;
	reg                r_sub06_U_r_w;
	wire signed [ 9:0] w_sub06_result_addr;
	reg  signed [ 9:0] r_sub06_result_addr;
	wire        [31:0] w_sub06_result_datain;
	reg         [31:0] r_sub06_result_datain;
	wire        [31:0] w_sub06_result_dataout;
	wire               w_sub06_result_r_w;
	reg                r_sub06_result_r_w;
	reg                r_sub05_run_req;
	wire               w_sub05_run_busy;
	wire signed [ 9:0] w_sub05_T_addr;
	reg  signed [ 9:0] r_sub05_T_addr;
	wire        [31:0] w_sub05_T_datain;
	reg         [31:0] r_sub05_T_datain;
	wire        [31:0] w_sub05_T_dataout;
	wire               w_sub05_T_r_w;
	reg                r_sub05_T_r_w;
	wire signed [ 9:0] w_sub05_V_addr;
	reg  signed [ 9:0] r_sub05_V_addr;
	wire        [31:0] w_sub05_V_datain;
	reg         [31:0] r_sub05_V_datain;
	wire        [31:0] w_sub05_V_dataout;
	wire               w_sub05_V_r_w;
	reg                r_sub05_V_r_w;
	wire signed [ 9:0] w_sub05_U_addr;
	reg  signed [ 9:0] r_sub05_U_addr;
	wire        [31:0] w_sub05_U_datain;
	reg         [31:0] r_sub05_U_datain;
	wire        [31:0] w_sub05_U_dataout;
	wire               w_sub05_U_r_w;
	reg                r_sub05_U_r_w;
	wire signed [ 9:0] w_sub05_result_addr;
	reg  signed [ 9:0] r_sub05_result_addr;
	wire        [31:0] w_sub05_result_datain;
	reg         [31:0] r_sub05_result_datain;
	wire        [31:0] w_sub05_result_dataout;
	wire               w_sub05_result_r_w;
	reg                r_sub05_result_r_w;
	reg                r_sub04_run_req;
	wire               w_sub04_run_busy;
	wire signed [ 9:0] w_sub04_T_addr;
	reg  signed [ 9:0] r_sub04_T_addr;
	wire        [31:0] w_sub04_T_datain;
	reg         [31:0] r_sub04_T_datain;
	wire        [31:0] w_sub04_T_dataout;
	wire               w_sub04_T_r_w;
	reg                r_sub04_T_r_w;
	wire signed [ 9:0] w_sub04_V_addr;
	reg  signed [ 9:0] r_sub04_V_addr;
	wire        [31:0] w_sub04_V_datain;
	reg         [31:0] r_sub04_V_datain;
	wire        [31:0] w_sub04_V_dataout;
	wire               w_sub04_V_r_w;
	reg                r_sub04_V_r_w;
	wire signed [ 9:0] w_sub04_U_addr;
	reg  signed [ 9:0] r_sub04_U_addr;
	wire        [31:0] w_sub04_U_datain;
	reg         [31:0] r_sub04_U_datain;
	wire        [31:0] w_sub04_U_dataout;
	wire               w_sub04_U_r_w;
	reg                r_sub04_U_r_w;
	wire signed [ 9:0] w_sub04_result_addr;
	reg  signed [ 9:0] r_sub04_result_addr;
	wire        [31:0] w_sub04_result_datain;
	reg         [31:0] r_sub04_result_datain;
	wire        [31:0] w_sub04_result_dataout;
	wire               w_sub04_result_r_w;
	reg                r_sub04_result_r_w;
	reg         [31:0] r_sys_tmp0_float;
	reg         [31:0] r_sys_tmp1_float;
	reg         [31:0] r_sys_tmp2_float;
	reg         [31:0] r_sys_tmp3_float;
	reg         [31:0] r_sys_tmp4_float;
	reg         [31:0] r_sys_tmp5_float;
	reg         [31:0] r_sys_tmp6_float;
	reg         [31:0] r_sys_tmp7_float;
	reg         [31:0] r_sys_tmp8_float;
	reg         [31:0] r_sys_tmp9_float;
	reg         [31:0] r_sys_tmp10_float;
	reg         [31:0] r_sys_tmp11_float;
	reg         [31:0] r_sys_tmp12_float;
	reg         [31:0] r_sys_tmp13_float;
	reg         [31:0] r_sys_tmp14_float;
	reg         [31:0] r_sys_tmp15_float;
	reg         [31:0] r_sys_tmp16_float;
	reg         [31:0] r_sys_tmp17_float;
	reg         [31:0] r_sys_tmp18_float;
	reg         [31:0] r_sys_tmp19_float;
	reg         [31:0] r_sys_tmp20_float;
	reg         [31:0] r_sys_tmp21_float;
	reg         [31:0] r_sys_tmp22_float;
	reg         [31:0] r_sys_tmp23_float;
	reg         [31:0] r_sys_tmp24_float;
	reg         [31:0] r_sys_tmp25_float;
	reg         [31:0] r_sys_tmp26_float;
	reg         [31:0] r_sys_tmp27_float;
	reg         [31:0] r_sys_tmp28_float;
	reg         [31:0] r_sys_tmp29_float;
	reg         [31:0] r_sys_tmp30_float;
	reg         [31:0] r_sys_tmp31_float;
	reg         [31:0] r_sys_tmp32_float;
	reg         [31:0] r_sys_tmp33_float;
	reg         [31:0] r_sys_tmp34_float;
	reg         [31:0] r_sys_tmp35_float;
	reg         [31:0] r_sys_tmp36_float;
	reg         [31:0] r_sys_tmp37_float;
	reg         [31:0] r_sys_tmp38_float;
	reg         [31:0] r_sys_tmp39_float;
	reg         [31:0] r_sys_tmp40_float;
	reg         [31:0] r_sys_tmp41_float;
	reg         [31:0] r_sys_tmp42_float;
	reg         [31:0] r_sys_tmp43_float;
	reg         [31:0] r_sys_tmp44_float;
	reg         [31:0] r_sys_tmp45_float;
	reg         [31:0] r_sys_tmp46_float;
	reg         [31:0] r_sys_tmp47_float;
	wire signed [31:0] w_sys_tmp1;
	wire signed [31:0] w_sys_tmp3;
	wire        [31:0] w_sys_tmp5;
	wire signed [31:0] w_sys_tmp6;
	wire        [31:0] w_sys_tmp7;
	wire        [31:0] w_sys_tmp8;
	wire        [31:0] w_sys_tmp9;
	wire        [31:0] w_sys_tmp10;
	wire        [31:0] w_sys_tmp11;
	wire        [31:0] w_sys_tmp12;
	wire               w_sys_tmp13;
	wire               w_sys_tmp14;
	wire signed [31:0] w_sys_tmp15;
	wire               w_sys_tmp16;
	wire               w_sys_tmp17;
	wire        [31:0] w_sys_tmp19;
	wire        [31:0] w_sys_tmp20;
	wire signed [31:0] w_sys_tmp21;
	wire signed [31:0] w_sys_tmp23;
	wire signed [31:0] w_sys_tmp24;
	wire signed [31:0] w_sys_tmp25;
	wire        [31:0] w_sys_tmp26;
	wire signed [31:0] w_sys_tmp28;
	wire signed [31:0] w_sys_tmp29;
	wire signed [31:0] w_sys_tmp33;
	wire signed [31:0] w_sys_tmp34;
	wire        [31:0] w_sys_tmp37;
	wire        [31:0] w_sys_tmp38;
	wire        [31:0] w_sys_tmp39;
	wire signed [31:0] w_sys_tmp42;
	wire signed [31:0] w_sys_tmp43;
	wire signed [31:0] w_sys_tmp46;
	wire signed [31:0] w_sys_tmp47;
	wire signed [31:0] w_sys_tmp48;
	wire signed [31:0] w_sys_tmp49;
	wire        [31:0] w_sys_tmp129;
	wire               w_sys_tmp227;
	wire               w_sys_tmp228;
	wire signed [31:0] w_sys_tmp229;
	wire signed [31:0] w_sys_tmp232;
	wire signed [31:0] w_sys_tmp233;
	wire        [31:0] w_sys_tmp234;
	wire        [31:0] w_sys_tmp240;
	wire signed [31:0] w_sys_tmp244;
	wire signed [31:0] w_sys_tmp245;
	wire signed [31:0] w_sys_tmp256;
	wire signed [31:0] w_sys_tmp257;
	wire signed [31:0] w_sys_tmp268;
	wire signed [31:0] w_sys_tmp269;
	wire signed [31:0] w_sys_tmp280;
	wire signed [31:0] w_sys_tmp281;
	wire signed [31:0] w_sys_tmp292;
	wire signed [31:0] w_sys_tmp293;
	wire signed [31:0] w_sys_tmp304;
	wire signed [31:0] w_sys_tmp305;
	wire signed [31:0] w_sys_tmp316;
	wire signed [31:0] w_sys_tmp317;
	wire signed [31:0] w_sys_tmp328;
	wire signed [31:0] w_sys_tmp329;
	wire signed [31:0] w_sys_tmp340;
	wire signed [31:0] w_sys_tmp341;
	wire signed [31:0] w_sys_tmp352;
	wire signed [31:0] w_sys_tmp353;
	wire signed [31:0] w_sys_tmp364;
	wire signed [31:0] w_sys_tmp365;
	wire signed [31:0] w_sys_tmp400;
	wire signed [31:0] w_sys_tmp401;
	wire signed [31:0] w_sys_tmp412;
	wire signed [31:0] w_sys_tmp413;
	wire signed [31:0] w_sys_tmp424;
	wire signed [31:0] w_sys_tmp425;
	wire signed [31:0] w_sys_tmp436;
	wire signed [31:0] w_sys_tmp437;
	wire signed [31:0] w_sys_tmp448;
	wire signed [31:0] w_sys_tmp449;
	wire signed [31:0] w_sys_tmp460;
	wire signed [31:0] w_sys_tmp461;
	wire signed [31:0] w_sys_tmp472;
	wire signed [31:0] w_sys_tmp473;
	wire signed [31:0] w_sys_tmp484;
	wire signed [31:0] w_sys_tmp485;
	wire signed [31:0] w_sys_tmp496;
	wire signed [31:0] w_sys_tmp497;
	wire signed [31:0] w_sys_tmp508;
	wire signed [31:0] w_sys_tmp509;
	wire signed [31:0] w_sys_tmp544;
	wire signed [31:0] w_sys_tmp545;
	wire signed [31:0] w_sys_tmp556;
	wire signed [31:0] w_sys_tmp557;
	wire signed [31:0] w_sys_tmp568;
	wire signed [31:0] w_sys_tmp569;
	wire signed [31:0] w_sys_tmp580;
	wire signed [31:0] w_sys_tmp581;
	wire signed [31:0] w_sys_tmp592;
	wire signed [31:0] w_sys_tmp593;
	wire signed [31:0] w_sys_tmp604;
	wire signed [31:0] w_sys_tmp605;
	wire signed [31:0] w_sys_tmp616;
	wire signed [31:0] w_sys_tmp617;
	wire signed [31:0] w_sys_tmp628;
	wire signed [31:0] w_sys_tmp629;
	wire signed [31:0] w_sys_tmp640;
	wire signed [31:0] w_sys_tmp641;
	wire signed [31:0] w_sys_tmp652;
	wire signed [31:0] w_sys_tmp653;
	wire signed [31:0] w_sys_tmp664;
	wire signed [31:0] w_sys_tmp665;
	wire signed [31:0] w_sys_tmp676;
	wire signed [31:0] w_sys_tmp677;
	wire signed [31:0] w_sys_tmp688;
	wire signed [31:0] w_sys_tmp689;
	wire signed [31:0] w_sys_tmp700;
	wire signed [31:0] w_sys_tmp701;
	wire signed [31:0] w_sys_tmp712;
	wire signed [31:0] w_sys_tmp713;
	wire signed [31:0] w_sys_tmp724;
	wire signed [31:0] w_sys_tmp725;
	wire signed [31:0] w_sys_tmp736;
	wire signed [31:0] w_sys_tmp737;
	wire signed [31:0] w_sys_tmp748;
	wire signed [31:0] w_sys_tmp749;
	wire signed [31:0] w_sys_tmp760;
	wire signed [31:0] w_sys_tmp761;
	wire signed [31:0] w_sys_tmp772;
	wire signed [31:0] w_sys_tmp773;
	wire signed [31:0] w_sys_tmp784;
	wire signed [31:0] w_sys_tmp785;
	wire signed [31:0] w_sys_tmp820;
	wire signed [31:0] w_sys_tmp821;
	wire signed [31:0] w_sys_tmp832;
	wire signed [31:0] w_sys_tmp833;
	wire signed [31:0] w_sys_tmp844;
	wire signed [31:0] w_sys_tmp845;
	wire signed [31:0] w_sys_tmp856;
	wire signed [31:0] w_sys_tmp857;
	wire signed [31:0] w_sys_tmp868;
	wire signed [31:0] w_sys_tmp869;
	wire signed [31:0] w_sys_tmp880;
	wire signed [31:0] w_sys_tmp881;
	wire signed [31:0] w_sys_tmp892;
	wire signed [31:0] w_sys_tmp893;
	wire signed [31:0] w_sys_tmp904;
	wire signed [31:0] w_sys_tmp905;
	wire signed [31:0] w_sys_tmp916;
	wire signed [31:0] w_sys_tmp917;
	wire signed [31:0] w_sys_tmp928;
	wire signed [31:0] w_sys_tmp929;
	wire signed [31:0] w_sys_tmp964;
	wire signed [31:0] w_sys_tmp965;
	wire signed [31:0] w_sys_tmp976;
	wire signed [31:0] w_sys_tmp977;
	wire signed [31:0] w_sys_tmp988;
	wire signed [31:0] w_sys_tmp989;
	wire signed [31:0] w_sys_tmp1000;
	wire signed [31:0] w_sys_tmp1001;
	wire signed [31:0] w_sys_tmp1012;
	wire signed [31:0] w_sys_tmp1013;
	wire signed [31:0] w_sys_tmp1024;
	wire signed [31:0] w_sys_tmp1025;
	wire signed [31:0] w_sys_tmp1036;
	wire signed [31:0] w_sys_tmp1037;
	wire signed [31:0] w_sys_tmp1048;
	wire signed [31:0] w_sys_tmp1049;
	wire signed [31:0] w_sys_tmp1060;
	wire signed [31:0] w_sys_tmp1061;
	wire signed [31:0] w_sys_tmp1071;
	wire signed [31:0] w_sys_tmp1072;
	wire               w_sys_tmp1073;
	wire               w_sys_tmp1074;
	wire signed [31:0] w_sys_tmp1075;
	wire signed [31:0] w_sys_tmp1078;
	wire signed [31:0] w_sys_tmp1079;
	wire        [31:0] w_sys_tmp1080;
	wire        [31:0] w_sys_tmp1086;
	wire signed [31:0] w_sys_tmp1090;
	wire signed [31:0] w_sys_tmp1091;
	wire signed [31:0] w_sys_tmp1102;
	wire signed [31:0] w_sys_tmp1103;
	wire signed [31:0] w_sys_tmp1114;
	wire signed [31:0] w_sys_tmp1115;
	wire signed [31:0] w_sys_tmp1126;
	wire signed [31:0] w_sys_tmp1127;
	wire signed [31:0] w_sys_tmp1138;
	wire signed [31:0] w_sys_tmp1139;
	wire signed [31:0] w_sys_tmp1150;
	wire signed [31:0] w_sys_tmp1151;
	wire signed [31:0] w_sys_tmp1162;
	wire signed [31:0] w_sys_tmp1163;
	wire signed [31:0] w_sys_tmp1174;
	wire signed [31:0] w_sys_tmp1175;
	wire signed [31:0] w_sys_tmp1186;
	wire signed [31:0] w_sys_tmp1187;
	wire signed [31:0] w_sys_tmp1198;
	wire signed [31:0] w_sys_tmp1199;
	wire signed [31:0] w_sys_tmp1210;
	wire signed [31:0] w_sys_tmp1211;
	wire signed [31:0] w_sys_tmp1246;
	wire signed [31:0] w_sys_tmp1247;
	wire signed [31:0] w_sys_tmp1258;
	wire signed [31:0] w_sys_tmp1259;
	wire signed [31:0] w_sys_tmp1270;
	wire signed [31:0] w_sys_tmp1271;
	wire signed [31:0] w_sys_tmp1282;
	wire signed [31:0] w_sys_tmp1283;
	wire signed [31:0] w_sys_tmp1294;
	wire signed [31:0] w_sys_tmp1295;
	wire signed [31:0] w_sys_tmp1306;
	wire signed [31:0] w_sys_tmp1307;
	wire signed [31:0] w_sys_tmp1318;
	wire signed [31:0] w_sys_tmp1319;
	wire signed [31:0] w_sys_tmp1330;
	wire signed [31:0] w_sys_tmp1331;
	wire signed [31:0] w_sys_tmp1342;
	wire signed [31:0] w_sys_tmp1343;
	wire signed [31:0] w_sys_tmp1366;
	wire signed [31:0] w_sys_tmp1367;
	wire signed [31:0] w_sys_tmp1378;
	wire signed [31:0] w_sys_tmp1379;
	wire signed [31:0] w_sys_tmp1390;
	wire signed [31:0] w_sys_tmp1391;
	wire signed [31:0] w_sys_tmp1402;
	wire signed [31:0] w_sys_tmp1403;
	wire signed [31:0] w_sys_tmp1414;
	wire signed [31:0] w_sys_tmp1415;
	wire signed [31:0] w_sys_tmp1426;
	wire signed [31:0] w_sys_tmp1427;
	wire signed [31:0] w_sys_tmp1438;
	wire signed [31:0] w_sys_tmp1439;
	wire signed [31:0] w_sys_tmp1450;
	wire signed [31:0] w_sys_tmp1451;
	wire signed [31:0] w_sys_tmp1462;
	wire signed [31:0] w_sys_tmp1463;
	wire signed [31:0] w_sys_tmp1473;
	wire               w_sys_tmp1474;
	wire               w_sys_tmp1475;
	wire signed [31:0] w_sys_tmp1476;
	wire               w_sys_tmp1477;
	wire               w_sys_tmp1478;
	wire signed [31:0] w_sys_tmp1481;
	wire signed [31:0] w_sys_tmp1482;
	wire        [31:0] w_sys_tmp1483;
	wire signed [31:0] w_sys_tmp1485;
	wire signed [31:0] w_sys_tmp1486;
	wire        [31:0] w_sys_tmp1488;
	wire signed [31:0] w_sys_tmp1489;
	wire signed [31:0] w_sys_tmp1490;
	wire signed [31:0] w_sys_tmp1491;
	wire signed [31:0] w_sys_tmp1493;
	wire               w_sys_tmp1494;
	wire               w_sys_tmp1495;
	wire signed [31:0] w_sys_tmp1498;
	wire signed [31:0] w_sys_tmp1499;
	wire signed [31:0] w_sys_tmp1500;
	wire        [31:0] w_sys_tmp1501;
	wire signed [31:0] w_sys_tmp1503;
	wire signed [31:0] w_sys_tmp1504;
	wire signed [31:0] w_sys_tmp1507;
	wire signed [31:0] w_sys_tmp1508;
	wire signed [31:0] w_sys_tmp1581;
	wire signed [31:0] w_sys_tmp1582;
	wire               w_sys_tmp1583;
	wire               w_sys_tmp1584;
	wire signed [31:0] w_sys_tmp1585;
	wire signed [31:0] w_sys_tmp1586;
	wire signed [31:0] w_sys_tmp1589;
	wire signed [31:0] w_sys_tmp1590;
	wire signed [31:0] w_sys_tmp1591;
	wire        [31:0] w_sys_tmp1592;
	wire signed [31:0] w_sys_tmp1593;
	wire               w_sys_tmp1630;
	wire               w_sys_tmp1631;
	wire signed [31:0] w_sys_tmp1632;
	wire signed [31:0] w_sys_tmp1635;
	wire signed [31:0] w_sys_tmp1636;
	wire        [31:0] w_sys_tmp1637;
	wire signed [31:0] w_sys_tmp1641;
	wire signed [31:0] w_sys_tmp1642;
	wire signed [31:0] w_sys_tmp1647;
	wire signed [31:0] w_sys_tmp1648;
	wire signed [31:0] w_sys_tmp1653;
	wire signed [31:0] w_sys_tmp1654;
	wire signed [31:0] w_sys_tmp1659;
	wire signed [31:0] w_sys_tmp1660;
	wire signed [31:0] w_sys_tmp1665;
	wire signed [31:0] w_sys_tmp1666;
	wire signed [31:0] w_sys_tmp1671;
	wire signed [31:0] w_sys_tmp1672;
	wire signed [31:0] w_sys_tmp1677;
	wire signed [31:0] w_sys_tmp1678;
	wire signed [31:0] w_sys_tmp1683;
	wire signed [31:0] w_sys_tmp1684;
	wire signed [31:0] w_sys_tmp1689;
	wire signed [31:0] w_sys_tmp1690;
	wire signed [31:0] w_sys_tmp1695;
	wire signed [31:0] w_sys_tmp1696;
	wire signed [31:0] w_sys_tmp1701;
	wire signed [31:0] w_sys_tmp1702;
	wire signed [31:0] w_sys_tmp1719;
	wire signed [31:0] w_sys_tmp1720;
	wire signed [31:0] w_sys_tmp1725;
	wire signed [31:0] w_sys_tmp1726;
	wire signed [31:0] w_sys_tmp1731;
	wire signed [31:0] w_sys_tmp1732;
	wire signed [31:0] w_sys_tmp1737;
	wire signed [31:0] w_sys_tmp1738;
	wire signed [31:0] w_sys_tmp1743;
	wire signed [31:0] w_sys_tmp1744;
	wire signed [31:0] w_sys_tmp1749;
	wire signed [31:0] w_sys_tmp1750;
	wire signed [31:0] w_sys_tmp1755;
	wire signed [31:0] w_sys_tmp1756;
	wire signed [31:0] w_sys_tmp1761;
	wire signed [31:0] w_sys_tmp1762;
	wire signed [31:0] w_sys_tmp1767;
	wire signed [31:0] w_sys_tmp1768;
	wire signed [31:0] w_sys_tmp1773;
	wire signed [31:0] w_sys_tmp1774;
	wire signed [31:0] w_sys_tmp1791;
	wire signed [31:0] w_sys_tmp1792;
	wire signed [31:0] w_sys_tmp1797;
	wire signed [31:0] w_sys_tmp1798;
	wire signed [31:0] w_sys_tmp1803;
	wire signed [31:0] w_sys_tmp1804;
	wire signed [31:0] w_sys_tmp1809;
	wire signed [31:0] w_sys_tmp1810;
	wire signed [31:0] w_sys_tmp1815;
	wire signed [31:0] w_sys_tmp1816;
	wire signed [31:0] w_sys_tmp1821;
	wire signed [31:0] w_sys_tmp1822;
	wire signed [31:0] w_sys_tmp1827;
	wire signed [31:0] w_sys_tmp1828;
	wire signed [31:0] w_sys_tmp1833;
	wire signed [31:0] w_sys_tmp1834;
	wire signed [31:0] w_sys_tmp1839;
	wire signed [31:0] w_sys_tmp1840;
	wire signed [31:0] w_sys_tmp1845;
	wire signed [31:0] w_sys_tmp1846;
	wire signed [31:0] w_sys_tmp1851;
	wire signed [31:0] w_sys_tmp1852;
	wire signed [31:0] w_sys_tmp1857;
	wire signed [31:0] w_sys_tmp1858;
	wire signed [31:0] w_sys_tmp1863;
	wire signed [31:0] w_sys_tmp1864;
	wire signed [31:0] w_sys_tmp1869;
	wire signed [31:0] w_sys_tmp1870;
	wire signed [31:0] w_sys_tmp1875;
	wire signed [31:0] w_sys_tmp1876;
	wire signed [31:0] w_sys_tmp1881;
	wire signed [31:0] w_sys_tmp1882;
	wire signed [31:0] w_sys_tmp1887;
	wire signed [31:0] w_sys_tmp1888;
	wire signed [31:0] w_sys_tmp1893;
	wire signed [31:0] w_sys_tmp1894;
	wire signed [31:0] w_sys_tmp1899;
	wire signed [31:0] w_sys_tmp1900;
	wire signed [31:0] w_sys_tmp1905;
	wire signed [31:0] w_sys_tmp1906;
	wire signed [31:0] w_sys_tmp1911;
	wire signed [31:0] w_sys_tmp1912;
	wire signed [31:0] w_sys_tmp1929;
	wire signed [31:0] w_sys_tmp1930;
	wire signed [31:0] w_sys_tmp1935;
	wire signed [31:0] w_sys_tmp1936;
	wire signed [31:0] w_sys_tmp1941;
	wire signed [31:0] w_sys_tmp1942;
	wire signed [31:0] w_sys_tmp1947;
	wire signed [31:0] w_sys_tmp1948;
	wire signed [31:0] w_sys_tmp1953;
	wire signed [31:0] w_sys_tmp1954;
	wire signed [31:0] w_sys_tmp1959;
	wire signed [31:0] w_sys_tmp1960;
	wire signed [31:0] w_sys_tmp1965;
	wire signed [31:0] w_sys_tmp1966;
	wire signed [31:0] w_sys_tmp1971;
	wire signed [31:0] w_sys_tmp1972;
	wire signed [31:0] w_sys_tmp1977;
	wire signed [31:0] w_sys_tmp1978;
	wire signed [31:0] w_sys_tmp1983;
	wire signed [31:0] w_sys_tmp1984;
	wire signed [31:0] w_sys_tmp2001;
	wire signed [31:0] w_sys_tmp2002;
	wire signed [31:0] w_sys_tmp2007;
	wire signed [31:0] w_sys_tmp2008;
	wire signed [31:0] w_sys_tmp2013;
	wire signed [31:0] w_sys_tmp2014;
	wire signed [31:0] w_sys_tmp2019;
	wire signed [31:0] w_sys_tmp2020;
	wire signed [31:0] w_sys_tmp2025;
	wire signed [31:0] w_sys_tmp2026;
	wire signed [31:0] w_sys_tmp2031;
	wire signed [31:0] w_sys_tmp2032;
	wire signed [31:0] w_sys_tmp2037;
	wire signed [31:0] w_sys_tmp2038;
	wire signed [31:0] w_sys_tmp2043;
	wire signed [31:0] w_sys_tmp2044;
	wire signed [31:0] w_sys_tmp2049;
	wire signed [31:0] w_sys_tmp2050;
	wire signed [31:0] w_sys_tmp2054;
	wire signed [31:0] w_sys_tmp2055;
	wire               w_sys_tmp2056;
	wire               w_sys_tmp2057;
	wire signed [31:0] w_sys_tmp2058;
	wire signed [31:0] w_sys_tmp2061;
	wire signed [31:0] w_sys_tmp2062;
	wire        [31:0] w_sys_tmp2063;
	wire signed [31:0] w_sys_tmp2067;
	wire signed [31:0] w_sys_tmp2068;
	wire signed [31:0] w_sys_tmp2073;
	wire signed [31:0] w_sys_tmp2074;
	wire signed [31:0] w_sys_tmp2079;
	wire signed [31:0] w_sys_tmp2080;
	wire signed [31:0] w_sys_tmp2085;
	wire signed [31:0] w_sys_tmp2086;
	wire signed [31:0] w_sys_tmp2091;
	wire signed [31:0] w_sys_tmp2092;
	wire signed [31:0] w_sys_tmp2097;
	wire signed [31:0] w_sys_tmp2098;
	wire signed [31:0] w_sys_tmp2103;
	wire signed [31:0] w_sys_tmp2104;
	wire signed [31:0] w_sys_tmp2109;
	wire signed [31:0] w_sys_tmp2110;
	wire signed [31:0] w_sys_tmp2115;
	wire signed [31:0] w_sys_tmp2116;
	wire signed [31:0] w_sys_tmp2121;
	wire signed [31:0] w_sys_tmp2122;
	wire signed [31:0] w_sys_tmp2127;
	wire signed [31:0] w_sys_tmp2128;
	wire signed [31:0] w_sys_tmp2145;
	wire signed [31:0] w_sys_tmp2146;
	wire signed [31:0] w_sys_tmp2151;
	wire signed [31:0] w_sys_tmp2152;
	wire signed [31:0] w_sys_tmp2157;
	wire signed [31:0] w_sys_tmp2158;
	wire signed [31:0] w_sys_tmp2163;
	wire signed [31:0] w_sys_tmp2164;
	wire signed [31:0] w_sys_tmp2169;
	wire signed [31:0] w_sys_tmp2170;
	wire signed [31:0] w_sys_tmp2175;
	wire signed [31:0] w_sys_tmp2176;
	wire signed [31:0] w_sys_tmp2181;
	wire signed [31:0] w_sys_tmp2182;
	wire signed [31:0] w_sys_tmp2187;
	wire signed [31:0] w_sys_tmp2188;
	wire signed [31:0] w_sys_tmp2193;
	wire signed [31:0] w_sys_tmp2194;
	wire signed [31:0] w_sys_tmp2199;
	wire signed [31:0] w_sys_tmp2200;
	wire signed [31:0] w_sys_tmp2217;
	wire signed [31:0] w_sys_tmp2218;
	wire signed [31:0] w_sys_tmp2223;
	wire signed [31:0] w_sys_tmp2224;
	wire signed [31:0] w_sys_tmp2229;
	wire signed [31:0] w_sys_tmp2230;
	wire signed [31:0] w_sys_tmp2235;
	wire signed [31:0] w_sys_tmp2236;
	wire signed [31:0] w_sys_tmp2241;
	wire signed [31:0] w_sys_tmp2242;
	wire signed [31:0] w_sys_tmp2247;
	wire signed [31:0] w_sys_tmp2248;
	wire signed [31:0] w_sys_tmp2253;
	wire signed [31:0] w_sys_tmp2254;
	wire signed [31:0] w_sys_tmp2259;
	wire signed [31:0] w_sys_tmp2260;
	wire signed [31:0] w_sys_tmp2264;
	wire signed [31:0] w_sys_tmp2265;
	wire               w_sys_tmp2266;
	wire               w_sys_tmp2267;
	wire signed [31:0] w_sys_tmp2268;
	wire signed [31:0] w_sys_tmp2271;
	wire signed [31:0] w_sys_tmp2272;
	wire        [31:0] w_sys_tmp2273;
	wire signed [31:0] w_sys_tmp2277;
	wire signed [31:0] w_sys_tmp2278;
	wire signed [31:0] w_sys_tmp2283;
	wire signed [31:0] w_sys_tmp2284;
	wire signed [31:0] w_sys_tmp2289;
	wire signed [31:0] w_sys_tmp2290;
	wire signed [31:0] w_sys_tmp2295;
	wire signed [31:0] w_sys_tmp2296;
	wire signed [31:0] w_sys_tmp2301;
	wire signed [31:0] w_sys_tmp2302;
	wire signed [31:0] w_sys_tmp2307;
	wire signed [31:0] w_sys_tmp2308;
	wire signed [31:0] w_sys_tmp2313;
	wire signed [31:0] w_sys_tmp2314;
	wire signed [31:0] w_sys_tmp2319;
	wire signed [31:0] w_sys_tmp2320;
	wire signed [31:0] w_sys_tmp2325;
	wire signed [31:0] w_sys_tmp2326;
	wire signed [31:0] w_sys_tmp2331;
	wire signed [31:0] w_sys_tmp2332;
	wire signed [31:0] w_sys_tmp2336;
	wire signed [31:0] w_sys_tmp2337;
	wire signed [31:0] w_sys_tmp2341;
	wire signed [31:0] w_sys_tmp2342;
	wire signed [31:0] w_sys_tmp2346;
	wire signed [31:0] w_sys_tmp2347;
	wire signed [31:0] w_sys_tmp2351;
	wire signed [31:0] w_sys_tmp2352;
	wire signed [31:0] w_sys_tmp2356;
	wire signed [31:0] w_sys_tmp2357;
	wire signed [31:0] w_sys_tmp2361;
	wire signed [31:0] w_sys_tmp2362;
	wire signed [31:0] w_sys_tmp2366;
	wire signed [31:0] w_sys_tmp2367;
	wire signed [31:0] w_sys_tmp2371;
	wire signed [31:0] w_sys_tmp2372;
	wire signed [31:0] w_sys_tmp2376;
	wire signed [31:0] w_sys_tmp2377;
	wire signed [31:0] w_sys_tmp2381;
	wire signed [31:0] w_sys_tmp2382;
	wire signed [31:0] w_sys_tmp2386;
	wire signed [31:0] w_sys_tmp2387;
	wire signed [31:0] w_sys_tmp2391;
	wire signed [31:0] w_sys_tmp2392;
	wire signed [31:0] w_sys_tmp2396;
	wire signed [31:0] w_sys_tmp2397;
	wire signed [31:0] w_sys_tmp2401;
	wire signed [31:0] w_sys_tmp2402;
	wire signed [31:0] w_sys_tmp2406;
	wire signed [31:0] w_sys_tmp2407;
	wire signed [31:0] w_sys_tmp2411;
	wire signed [31:0] w_sys_tmp2412;
	wire signed [31:0] w_sys_tmp2416;
	wire signed [31:0] w_sys_tmp2417;
	wire signed [31:0] w_sys_tmp2421;
	wire signed [31:0] w_sys_tmp2422;
	wire signed [31:0] w_sys_tmp2426;
	wire signed [31:0] w_sys_tmp2427;
	wire signed [31:0] w_sys_tmp2431;
	wire signed [31:0] w_sys_tmp2432;
	wire signed [31:0] w_sys_tmp2436;
	wire signed [31:0] w_sys_tmp2437;
	wire signed [31:0] w_sys_tmp2441;
	wire signed [31:0] w_sys_tmp2442;
	wire signed [31:0] w_sys_tmp2446;
	wire signed [31:0] w_sys_tmp2447;
	wire signed [31:0] w_sys_tmp2451;
	wire signed [31:0] w_sys_tmp2452;
	wire signed [31:0] w_sys_tmp2456;
	wire signed [31:0] w_sys_tmp2457;
	wire signed [31:0] w_sys_tmp2461;
	wire signed [31:0] w_sys_tmp2462;
	wire signed [31:0] w_sys_tmp2466;
	wire signed [31:0] w_sys_tmp2467;
	wire signed [31:0] w_sys_tmp2471;
	wire signed [31:0] w_sys_tmp2472;
	wire signed [31:0] w_sys_tmp2476;
	wire signed [31:0] w_sys_tmp2477;
	wire signed [31:0] w_sys_tmp2481;
	wire signed [31:0] w_sys_tmp2482;
	wire signed [31:0] w_sys_tmp2486;
	wire signed [31:0] w_sys_tmp2487;
	wire signed [31:0] w_sys_tmp2491;
	wire signed [31:0] w_sys_tmp2492;
	wire signed [31:0] w_sys_tmp2496;
	wire signed [31:0] w_sys_tmp2497;
	wire signed [31:0] w_sys_tmp2501;
	wire signed [31:0] w_sys_tmp2502;
	wire signed [31:0] w_sys_tmp2506;
	wire signed [31:0] w_sys_tmp2507;
	wire signed [31:0] w_sys_tmp2511;
	wire signed [31:0] w_sys_tmp2512;
	wire signed [31:0] w_sys_tmp2516;
	wire signed [31:0] w_sys_tmp2517;
	wire signed [31:0] w_sys_tmp2521;
	wire signed [31:0] w_sys_tmp2522;
	wire signed [31:0] w_sys_tmp2526;
	wire signed [31:0] w_sys_tmp2527;
	wire signed [31:0] w_sys_tmp2531;
	wire signed [31:0] w_sys_tmp2532;
	wire signed [31:0] w_sys_tmp2536;
	wire signed [31:0] w_sys_tmp2537;
	wire signed [31:0] w_sys_tmp2541;
	wire signed [31:0] w_sys_tmp2542;
	wire signed [31:0] w_sys_tmp2546;
	wire signed [31:0] w_sys_tmp2547;
	wire signed [31:0] w_sys_tmp2551;
	wire signed [31:0] w_sys_tmp2552;
	wire signed [31:0] w_sys_tmp2556;
	wire signed [31:0] w_sys_tmp2557;
	wire signed [31:0] w_sys_tmp2561;
	wire signed [31:0] w_sys_tmp2562;
	wire signed [31:0] w_sys_tmp2566;
	wire signed [31:0] w_sys_tmp2567;
	wire signed [31:0] w_sys_tmp2570;
	wire signed [31:0] w_sys_tmp2571;
	wire               w_sys_tmp2572;
	wire               w_sys_tmp2573;
	wire signed [31:0] w_sys_tmp2574;
	wire signed [31:0] w_sys_tmp2577;
	wire signed [31:0] w_sys_tmp2578;
	wire        [31:0] w_sys_tmp2579;
	wire signed [31:0] w_sys_tmp2583;
	wire signed [31:0] w_sys_tmp2584;
	wire signed [31:0] w_sys_tmp2589;
	wire signed [31:0] w_sys_tmp2590;
	wire signed [31:0] w_sys_tmp2595;
	wire signed [31:0] w_sys_tmp2596;
	wire signed [31:0] w_sys_tmp2601;
	wire signed [31:0] w_sys_tmp2602;
	wire signed [31:0] w_sys_tmp2607;
	wire signed [31:0] w_sys_tmp2608;
	wire signed [31:0] w_sys_tmp2613;
	wire signed [31:0] w_sys_tmp2614;
	wire signed [31:0] w_sys_tmp2619;
	wire signed [31:0] w_sys_tmp2620;
	wire signed [31:0] w_sys_tmp2625;
	wire signed [31:0] w_sys_tmp2626;
	wire signed [31:0] w_sys_tmp2631;
	wire signed [31:0] w_sys_tmp2632;
	wire signed [31:0] w_sys_tmp2637;
	wire signed [31:0] w_sys_tmp2638;
	wire signed [31:0] w_sys_tmp2642;
	wire signed [31:0] w_sys_tmp2643;
	wire signed [31:0] w_sys_tmp2647;
	wire signed [31:0] w_sys_tmp2648;
	wire signed [31:0] w_sys_tmp2652;
	wire signed [31:0] w_sys_tmp2653;
	wire signed [31:0] w_sys_tmp2657;
	wire signed [31:0] w_sys_tmp2658;
	wire signed [31:0] w_sys_tmp2662;
	wire signed [31:0] w_sys_tmp2663;
	wire signed [31:0] w_sys_tmp2667;
	wire signed [31:0] w_sys_tmp2668;
	wire signed [31:0] w_sys_tmp2672;
	wire signed [31:0] w_sys_tmp2673;
	wire signed [31:0] w_sys_tmp2677;
	wire signed [31:0] w_sys_tmp2678;
	wire signed [31:0] w_sys_tmp2682;
	wire signed [31:0] w_sys_tmp2683;
	wire signed [31:0] w_sys_tmp2687;
	wire signed [31:0] w_sys_tmp2688;
	wire signed [31:0] w_sys_tmp2692;
	wire signed [31:0] w_sys_tmp2693;
	wire signed [31:0] w_sys_tmp2697;
	wire signed [31:0] w_sys_tmp2698;
	wire signed [31:0] w_sys_tmp2702;
	wire signed [31:0] w_sys_tmp2703;
	wire signed [31:0] w_sys_tmp2707;
	wire signed [31:0] w_sys_tmp2708;
	wire signed [31:0] w_sys_tmp2712;
	wire signed [31:0] w_sys_tmp2713;
	wire signed [31:0] w_sys_tmp2717;
	wire signed [31:0] w_sys_tmp2718;
	wire signed [31:0] w_sys_tmp2722;
	wire signed [31:0] w_sys_tmp2723;
	wire signed [31:0] w_sys_tmp2727;
	wire signed [31:0] w_sys_tmp2728;
	wire signed [31:0] w_sys_tmp2731;

	assign w_sys_boolTrue = 1'b1;
	assign w_sys_boolFalse = 1'b0;
	assign w_sys_intOne = 32'sh1;
	assign w_sys_intZero = 32'sh0;
	assign w_sys_ce = w_sys_boolTrue & ce;
	assign o_run_busy = r_sys_run_busy;
	assign w_sys_run_stage_p1 = (r_sys_run_stage + 4'h1);
	assign w_sys_run_step_p1 = (r_sys_run_step + 7'h1);
	assign w_fld_T_0_addr_0 = 9'sh0;
	assign w_fld_T_0_datain_0 = 32'h0;
	assign w_fld_T_0_r_w_0 = 1'h0;
	assign w_fld_T_0_ce_0 = w_sys_ce;
	assign w_fld_T_0_ce_1 = w_sys_ce;
	assign w_fld_TT_1_addr_0 = 9'sh0;
	assign w_fld_TT_1_datain_0 = 32'h0;
	assign w_fld_TT_1_r_w_0 = 1'h0;
	assign w_fld_TT_1_ce_0 = w_sys_ce;
	assign w_fld_TT_1_ce_1 = w_sys_ce;
	assign w_fld_U_2_addr_0 = 9'sh0;
	assign w_fld_U_2_datain_0 = 32'h0;
	assign w_fld_U_2_r_w_0 = 1'h0;
	assign w_fld_U_2_ce_0 = w_sys_ce;
	assign w_fld_U_2_ce_1 = w_sys_ce;
	assign w_fld_V_3_addr_0 = 9'sh0;
	assign w_fld_V_3_datain_0 = 32'h0;
	assign w_fld_V_3_r_w_0 = 1'h0;
	assign w_fld_V_3_ce_0 = w_sys_ce;
	assign w_fld_V_3_ce_1 = w_sys_ce;
	assign w_sub08_T_addr = ( (|r_sys_processing_methodID) ? r_sub08_T_addr : 10'sh0 ) ;
	assign w_sub08_T_datain = ( (|r_sys_processing_methodID) ? r_sub08_T_datain : 32'h0 ) ;
	assign w_sub08_T_r_w = ( (|r_sys_processing_methodID) ? r_sub08_T_r_w : 1'h0 ) ;
	assign w_sub08_V_addr = ( (|r_sys_processing_methodID) ? r_sub08_V_addr : 10'sh0 ) ;
	assign w_sub08_V_datain = ( (|r_sys_processing_methodID) ? r_sub08_V_datain : 32'h0 ) ;
	assign w_sub08_V_r_w = ( (|r_sys_processing_methodID) ? r_sub08_V_r_w : 1'h0 ) ;
	assign w_sub08_U_addr = ( (|r_sys_processing_methodID) ? r_sub08_U_addr : 10'sh0 ) ;
	assign w_sub08_U_datain = ( (|r_sys_processing_methodID) ? r_sub08_U_datain : 32'h0 ) ;
	assign w_sub08_U_r_w = ( (|r_sys_processing_methodID) ? r_sub08_U_r_w : 1'h0 ) ;
	assign w_sub08_result_addr = ( (|r_sys_processing_methodID) ? r_sub08_result_addr : 10'sh0 ) ;
	assign w_sub08_result_datain = ( (|r_sys_processing_methodID) ? r_sub08_result_datain : 32'h0 ) ;
	assign w_sub08_result_r_w = ( (|r_sys_processing_methodID) ? r_sub08_result_r_w : 1'h0 ) ;
	assign w_sub03_T_addr = ( (|r_sys_processing_methodID) ? r_sub03_T_addr : 10'sh0 ) ;
	assign w_sub03_T_datain = ( (|r_sys_processing_methodID) ? r_sub03_T_datain : 32'h0 ) ;
	assign w_sub03_T_r_w = ( (|r_sys_processing_methodID) ? r_sub03_T_r_w : 1'h0 ) ;
	assign w_sub03_V_addr = ( (|r_sys_processing_methodID) ? r_sub03_V_addr : 10'sh0 ) ;
	assign w_sub03_V_datain = ( (|r_sys_processing_methodID) ? r_sub03_V_datain : 32'h0 ) ;
	assign w_sub03_V_r_w = ( (|r_sys_processing_methodID) ? r_sub03_V_r_w : 1'h0 ) ;
	assign w_sub03_U_addr = ( (|r_sys_processing_methodID) ? r_sub03_U_addr : 10'sh0 ) ;
	assign w_sub03_U_datain = ( (|r_sys_processing_methodID) ? r_sub03_U_datain : 32'h0 ) ;
	assign w_sub03_U_r_w = ( (|r_sys_processing_methodID) ? r_sub03_U_r_w : 1'h0 ) ;
	assign w_sub03_result_addr = ( (|r_sys_processing_methodID) ? r_sub03_result_addr : 10'sh0 ) ;
	assign w_sub03_result_datain = ( (|r_sys_processing_methodID) ? r_sub03_result_datain : 32'h0 ) ;
	assign w_sub03_result_r_w = ( (|r_sys_processing_methodID) ? r_sub03_result_r_w : 1'h0 ) ;
	assign w_sub02_T_addr = ( (|r_sys_processing_methodID) ? r_sub02_T_addr : 10'sh0 ) ;
	assign w_sub02_T_datain = ( (|r_sys_processing_methodID) ? r_sub02_T_datain : 32'h0 ) ;
	assign w_sub02_T_r_w = ( (|r_sys_processing_methodID) ? r_sub02_T_r_w : 1'h0 ) ;
	assign w_sub02_V_addr = ( (|r_sys_processing_methodID) ? r_sub02_V_addr : 10'sh0 ) ;
	assign w_sub02_V_datain = ( (|r_sys_processing_methodID) ? r_sub02_V_datain : 32'h0 ) ;
	assign w_sub02_V_r_w = ( (|r_sys_processing_methodID) ? r_sub02_V_r_w : 1'h0 ) ;
	assign w_sub02_U_addr = ( (|r_sys_processing_methodID) ? r_sub02_U_addr : 10'sh0 ) ;
	assign w_sub02_U_datain = ( (|r_sys_processing_methodID) ? r_sub02_U_datain : 32'h0 ) ;
	assign w_sub02_U_r_w = ( (|r_sys_processing_methodID) ? r_sub02_U_r_w : 1'h0 ) ;
	assign w_sub02_result_addr = ( (|r_sys_processing_methodID) ? r_sub02_result_addr : 10'sh0 ) ;
	assign w_sub02_result_datain = ( (|r_sys_processing_methodID) ? r_sub02_result_datain : 32'h0 ) ;
	assign w_sub02_result_r_w = ( (|r_sys_processing_methodID) ? r_sub02_result_r_w : 1'h0 ) ;
	assign w_sub01_T_addr = ( (|r_sys_processing_methodID) ? r_sub01_T_addr : 10'sh0 ) ;
	assign w_sub01_T_datain = ( (|r_sys_processing_methodID) ? r_sub01_T_datain : 32'h0 ) ;
	assign w_sub01_T_r_w = ( (|r_sys_processing_methodID) ? r_sub01_T_r_w : 1'h0 ) ;
	assign w_sub01_V_addr = ( (|r_sys_processing_methodID) ? r_sub01_V_addr : 10'sh0 ) ;
	assign w_sub01_V_datain = ( (|r_sys_processing_methodID) ? r_sub01_V_datain : 32'h0 ) ;
	assign w_sub01_V_r_w = ( (|r_sys_processing_methodID) ? r_sub01_V_r_w : 1'h0 ) ;
	assign w_sub01_U_addr = ( (|r_sys_processing_methodID) ? r_sub01_U_addr : 10'sh0 ) ;
	assign w_sub01_U_datain = ( (|r_sys_processing_methodID) ? r_sub01_U_datain : 32'h0 ) ;
	assign w_sub01_U_r_w = ( (|r_sys_processing_methodID) ? r_sub01_U_r_w : 1'h0 ) ;
	assign w_sub01_result_addr = ( (|r_sys_processing_methodID) ? r_sub01_result_addr : 10'sh0 ) ;
	assign w_sub01_result_datain = ( (|r_sys_processing_methodID) ? r_sub01_result_datain : 32'h0 ) ;
	assign w_sub01_result_r_w = ( (|r_sys_processing_methodID) ? r_sub01_result_r_w : 1'h0 ) ;
	assign w_sub00_T_addr = ( (|r_sys_processing_methodID) ? r_sub00_T_addr : 10'sh0 ) ;
	assign w_sub00_T_datain = ( (|r_sys_processing_methodID) ? r_sub00_T_datain : 32'h0 ) ;
	assign w_sub00_T_r_w = ( (|r_sys_processing_methodID) ? r_sub00_T_r_w : 1'h0 ) ;
	assign w_sub00_V_addr = ( (|r_sys_processing_methodID) ? r_sub00_V_addr : 10'sh0 ) ;
	assign w_sub00_V_datain = ( (|r_sys_processing_methodID) ? r_sub00_V_datain : 32'h0 ) ;
	assign w_sub00_V_r_w = ( (|r_sys_processing_methodID) ? r_sub00_V_r_w : 1'h0 ) ;
	assign w_sub00_U_addr = ( (|r_sys_processing_methodID) ? r_sub00_U_addr : 10'sh0 ) ;
	assign w_sub00_U_datain = ( (|r_sys_processing_methodID) ? r_sub00_U_datain : 32'h0 ) ;
	assign w_sub00_U_r_w = ( (|r_sys_processing_methodID) ? r_sub00_U_r_w : 1'h0 ) ;
	assign w_sub00_result_addr = ( (|r_sys_processing_methodID) ? r_sub00_result_addr : 10'sh0 ) ;
	assign w_sub00_result_datain = ( (|r_sys_processing_methodID) ? r_sub00_result_datain : 32'h0 ) ;
	assign w_sub00_result_r_w = ( (|r_sys_processing_methodID) ? r_sub00_result_r_w : 1'h0 ) ;
	assign w_sub07_T_addr = ( (|r_sys_processing_methodID) ? r_sub07_T_addr : 10'sh0 ) ;
	assign w_sub07_T_datain = ( (|r_sys_processing_methodID) ? r_sub07_T_datain : 32'h0 ) ;
	assign w_sub07_T_r_w = ( (|r_sys_processing_methodID) ? r_sub07_T_r_w : 1'h0 ) ;
	assign w_sub07_V_addr = ( (|r_sys_processing_methodID) ? r_sub07_V_addr : 10'sh0 ) ;
	assign w_sub07_V_datain = ( (|r_sys_processing_methodID) ? r_sub07_V_datain : 32'h0 ) ;
	assign w_sub07_V_r_w = ( (|r_sys_processing_methodID) ? r_sub07_V_r_w : 1'h0 ) ;
	assign w_sub07_U_addr = ( (|r_sys_processing_methodID) ? r_sub07_U_addr : 10'sh0 ) ;
	assign w_sub07_U_datain = ( (|r_sys_processing_methodID) ? r_sub07_U_datain : 32'h0 ) ;
	assign w_sub07_U_r_w = ( (|r_sys_processing_methodID) ? r_sub07_U_r_w : 1'h0 ) ;
	assign w_sub07_result_addr = ( (|r_sys_processing_methodID) ? r_sub07_result_addr : 10'sh0 ) ;
	assign w_sub07_result_datain = ( (|r_sys_processing_methodID) ? r_sub07_result_datain : 32'h0 ) ;
	assign w_sub07_result_r_w = ( (|r_sys_processing_methodID) ? r_sub07_result_r_w : 1'h0 ) ;
	assign w_sub06_T_addr = ( (|r_sys_processing_methodID) ? r_sub06_T_addr : 10'sh0 ) ;
	assign w_sub06_T_datain = ( (|r_sys_processing_methodID) ? r_sub06_T_datain : 32'h0 ) ;
	assign w_sub06_T_r_w = ( (|r_sys_processing_methodID) ? r_sub06_T_r_w : 1'h0 ) ;
	assign w_sub06_V_addr = ( (|r_sys_processing_methodID) ? r_sub06_V_addr : 10'sh0 ) ;
	assign w_sub06_V_datain = ( (|r_sys_processing_methodID) ? r_sub06_V_datain : 32'h0 ) ;
	assign w_sub06_V_r_w = ( (|r_sys_processing_methodID) ? r_sub06_V_r_w : 1'h0 ) ;
	assign w_sub06_U_addr = ( (|r_sys_processing_methodID) ? r_sub06_U_addr : 10'sh0 ) ;
	assign w_sub06_U_datain = ( (|r_sys_processing_methodID) ? r_sub06_U_datain : 32'h0 ) ;
	assign w_sub06_U_r_w = ( (|r_sys_processing_methodID) ? r_sub06_U_r_w : 1'h0 ) ;
	assign w_sub06_result_addr = ( (|r_sys_processing_methodID) ? r_sub06_result_addr : 10'sh0 ) ;
	assign w_sub06_result_datain = ( (|r_sys_processing_methodID) ? r_sub06_result_datain : 32'h0 ) ;
	assign w_sub06_result_r_w = ( (|r_sys_processing_methodID) ? r_sub06_result_r_w : 1'h0 ) ;
	assign w_sub05_T_addr = ( (|r_sys_processing_methodID) ? r_sub05_T_addr : 10'sh0 ) ;
	assign w_sub05_T_datain = ( (|r_sys_processing_methodID) ? r_sub05_T_datain : 32'h0 ) ;
	assign w_sub05_T_r_w = ( (|r_sys_processing_methodID) ? r_sub05_T_r_w : 1'h0 ) ;
	assign w_sub05_V_addr = ( (|r_sys_processing_methodID) ? r_sub05_V_addr : 10'sh0 ) ;
	assign w_sub05_V_datain = ( (|r_sys_processing_methodID) ? r_sub05_V_datain : 32'h0 ) ;
	assign w_sub05_V_r_w = ( (|r_sys_processing_methodID) ? r_sub05_V_r_w : 1'h0 ) ;
	assign w_sub05_U_addr = ( (|r_sys_processing_methodID) ? r_sub05_U_addr : 10'sh0 ) ;
	assign w_sub05_U_datain = ( (|r_sys_processing_methodID) ? r_sub05_U_datain : 32'h0 ) ;
	assign w_sub05_U_r_w = ( (|r_sys_processing_methodID) ? r_sub05_U_r_w : 1'h0 ) ;
	assign w_sub05_result_addr = ( (|r_sys_processing_methodID) ? r_sub05_result_addr : 10'sh0 ) ;
	assign w_sub05_result_datain = ( (|r_sys_processing_methodID) ? r_sub05_result_datain : 32'h0 ) ;
	assign w_sub05_result_r_w = ( (|r_sys_processing_methodID) ? r_sub05_result_r_w : 1'h0 ) ;
	assign w_sub04_T_addr = ( (|r_sys_processing_methodID) ? r_sub04_T_addr : 10'sh0 ) ;
	assign w_sub04_T_datain = ( (|r_sys_processing_methodID) ? r_sub04_T_datain : 32'h0 ) ;
	assign w_sub04_T_r_w = ( (|r_sys_processing_methodID) ? r_sub04_T_r_w : 1'h0 ) ;
	assign w_sub04_V_addr = ( (|r_sys_processing_methodID) ? r_sub04_V_addr : 10'sh0 ) ;
	assign w_sub04_V_datain = ( (|r_sys_processing_methodID) ? r_sub04_V_datain : 32'h0 ) ;
	assign w_sub04_V_r_w = ( (|r_sys_processing_methodID) ? r_sub04_V_r_w : 1'h0 ) ;
	assign w_sub04_U_addr = ( (|r_sys_processing_methodID) ? r_sub04_U_addr : 10'sh0 ) ;
	assign w_sub04_U_datain = ( (|r_sys_processing_methodID) ? r_sub04_U_datain : 32'h0 ) ;
	assign w_sub04_U_r_w = ( (|r_sys_processing_methodID) ? r_sub04_U_r_w : 1'h0 ) ;
	assign w_sub04_result_addr = ( (|r_sys_processing_methodID) ? r_sub04_result_addr : 10'sh0 ) ;
	assign w_sub04_result_datain = ( (|r_sys_processing_methodID) ? r_sub04_result_datain : 32'h0 ) ;
	assign w_sub04_result_r_w = ( (|r_sys_processing_methodID) ? r_sub04_result_r_w : 1'h0 ) ;
	assign w_sys_tmp1 = 32'sh0000001e;
	assign w_sys_tmp3 = 32'sh0000001f;
	assign w_sys_tmp5 = 32'h3a03126f;
	assign w_sys_tmp6 = 32'sh00000190;
	assign w_sys_tmp7 = 32'h3e088889;
	assign w_sys_tmp8 = 32'h3d088889;
	assign w_sys_tmp9 = 32'h3af5c28f;
	assign w_sys_tmp10 = 32'h3bf5c28f;
	assign w_sys_tmp11 = 32'h3ce66665;
	assign w_sys_tmp12 = 32'h3ee66665;
	assign w_sys_tmp13 = ( !w_sys_tmp14 );
	assign w_sys_tmp14 = (r_run_my_17 < r_run_k_13);
	assign w_sys_tmp15 = (r_run_k_13 + w_sys_intOne);
	assign w_sys_tmp16 = ( !w_sys_tmp17 );
	assign w_sys_tmp17 = (r_run_mx_16 < r_run_j_14);
	assign w_sys_tmp19 = w_ip_MultFloat_product_0;
	assign w_sys_tmp20 = w_ip_FixedToFloat_floating_0;
	assign w_sys_tmp21 = (r_run_k_13 - w_sys_intOne);
	assign w_sys_tmp23 = (w_sys_tmp24 + r_run_k_13);
	assign w_sys_tmp24 = (r_run_j_14 * w_sys_tmp25);
	assign w_sys_tmp25 = 32'sh0000001f;
	assign w_sys_tmp26 = 32'h0;
	assign w_sys_tmp28 = (w_sys_tmp29 + r_run_k_13);
	assign w_sys_tmp29 = (r_run_copy2_j_31 * w_sys_tmp25);
	assign w_sys_tmp33 = (w_sys_tmp34 + r_run_k_13);
	assign w_sys_tmp34 = (r_run_copy1_j_30 * w_sys_tmp25);
	assign w_sys_tmp37 = 32'h42200000;
	assign w_sys_tmp38 = w_sys_tmp19;
	assign w_sys_tmp39 = 32'h3f800000;
	assign w_sys_tmp42 = (w_sys_tmp43 + r_run_k_13);
	assign w_sys_tmp43 = (r_run_copy0_j_29 * w_sys_tmp25);
	assign w_sys_tmp46 = (r_run_copy0_j_29 + w_sys_intOne);
	assign w_sys_tmp47 = (r_run_copy1_j_30 + w_sys_intOne);
	assign w_sys_tmp48 = (r_run_copy2_j_31 + w_sys_intOne);
	assign w_sys_tmp49 = (r_run_j_14 + w_sys_intOne);
	assign w_sys_tmp129 = r_sys_tmp4_float;
	assign w_sys_tmp227 = ( !w_sys_tmp228 );
	assign w_sys_tmp228 = (w_sys_tmp229 < r_run_k_13);
	assign w_sys_tmp229 = 32'sh0000000c;
	assign w_sys_tmp232 = (w_sys_tmp233 + r_run_k_13);
	assign w_sys_tmp233 = 32'sh0000001f;
	assign w_sys_tmp234 = w_fld_U_2_dataout_1;
	assign w_sys_tmp240 = w_fld_V_3_dataout_1;
	assign w_sys_tmp244 = (w_sys_tmp245 + r_run_k_13);
	assign w_sys_tmp245 = 32'sh0000003e;
	assign w_sys_tmp256 = (w_sys_tmp257 + r_run_k_13);
	assign w_sys_tmp257 = 32'sh0000005d;
	assign w_sys_tmp268 = (w_sys_tmp269 + r_run_k_13);
	assign w_sys_tmp269 = 32'sh0000007c;
	assign w_sys_tmp280 = (w_sys_tmp281 + r_run_k_13);
	assign w_sys_tmp281 = 32'sh0000009b;
	assign w_sys_tmp292 = (w_sys_tmp293 + r_run_k_13);
	assign w_sys_tmp293 = 32'sh000000ba;
	assign w_sys_tmp304 = (w_sys_tmp305 + r_run_k_13);
	assign w_sys_tmp305 = 32'sh000000d9;
	assign w_sys_tmp316 = (w_sys_tmp317 + r_run_k_13);
	assign w_sys_tmp317 = 32'sh000000f8;
	assign w_sys_tmp328 = (w_sys_tmp329 + r_run_k_13);
	assign w_sys_tmp329 = 32'sh00000117;
	assign w_sys_tmp340 = (w_sys_tmp341 + r_run_k_13);
	assign w_sys_tmp341 = 32'sh00000136;
	assign w_sys_tmp352 = (w_sys_tmp353 + r_run_k_13);
	assign w_sys_tmp353 = 32'sh00000155;
	assign w_sys_tmp364 = (w_sys_tmp365 + r_run_k_13);
	assign w_sys_tmp365 = 32'sh00000174;
	assign w_sys_tmp400 = (w_sys_tmp401 + r_run_k_13);
	assign w_sys_tmp401 = 32'sh00000193;
	assign w_sys_tmp412 = (w_sys_tmp413 + r_run_k_13);
	assign w_sys_tmp413 = 32'sh000001b2;
	assign w_sys_tmp424 = (w_sys_tmp425 + r_run_k_13);
	assign w_sys_tmp425 = 32'sh000001d1;
	assign w_sys_tmp436 = (w_sys_tmp437 + r_run_k_13);
	assign w_sys_tmp437 = 32'sh000001f0;
	assign w_sys_tmp448 = (w_sys_tmp449 + r_run_k_13);
	assign w_sys_tmp449 = 32'sh0000020f;
	assign w_sys_tmp460 = (w_sys_tmp461 + r_run_k_13);
	assign w_sys_tmp461 = 32'sh0000022e;
	assign w_sys_tmp472 = (w_sys_tmp473 + r_run_k_13);
	assign w_sys_tmp473 = 32'sh0000024d;
	assign w_sys_tmp484 = (w_sys_tmp485 + r_run_k_13);
	assign w_sys_tmp485 = 32'sh0000026c;
	assign w_sys_tmp496 = (w_sys_tmp497 + r_run_k_13);
	assign w_sys_tmp497 = 32'sh0000028b;
	assign w_sys_tmp508 = (w_sys_tmp509 + r_run_k_13);
	assign w_sys_tmp509 = 32'sh000002aa;
	assign w_sys_tmp544 = (w_sys_tmp545 + r_run_k_13);
	assign w_sys_tmp545 = 32'sh000002c9;
	assign w_sys_tmp556 = (w_sys_tmp557 + r_run_k_13);
	assign w_sys_tmp557 = 32'sh000002e8;
	assign w_sys_tmp568 = (w_sys_tmp569 + r_run_k_13);
	assign w_sys_tmp569 = 32'sh00000307;
	assign w_sys_tmp580 = (w_sys_tmp581 + r_run_k_13);
	assign w_sys_tmp581 = 32'sh00000326;
	assign w_sys_tmp592 = (w_sys_tmp593 + r_run_k_13);
	assign w_sys_tmp593 = 32'sh00000345;
	assign w_sys_tmp604 = (w_sys_tmp605 + r_run_k_13);
	assign w_sys_tmp605 = 32'sh00000364;
	assign w_sys_tmp616 = (w_sys_tmp617 + r_run_k_13);
	assign w_sys_tmp617 = 32'sh00000383;
	assign w_sys_tmp628 = (w_sys_tmp629 + r_run_k_13);
	assign w_sys_tmp629 = 32'sh000003a2;
	assign w_sys_tmp640 = (w_sys_tmp641 + r_run_k_13);
	assign w_sys_tmp641 = 32'sh000003c1;
	assign w_sys_tmp652 = (w_sys_tmp653 + r_run_k_13);
	assign w_sys_tmp653 = 32'sh00000029;
	assign w_sys_tmp664 = (w_sys_tmp665 + r_run_k_13);
	assign w_sys_tmp665 = 32'sh00000048;
	assign w_sys_tmp676 = (w_sys_tmp677 + r_run_k_13);
	assign w_sys_tmp677 = 32'sh00000067;
	assign w_sys_tmp688 = (w_sys_tmp689 + r_run_k_13);
	assign w_sys_tmp689 = 32'sh00000086;
	assign w_sys_tmp700 = (w_sys_tmp701 + r_run_k_13);
	assign w_sys_tmp701 = 32'sh000000a5;
	assign w_sys_tmp712 = (w_sys_tmp713 + r_run_k_13);
	assign w_sys_tmp713 = 32'sh000000c4;
	assign w_sys_tmp724 = (w_sys_tmp725 + r_run_k_13);
	assign w_sys_tmp725 = 32'sh000000e3;
	assign w_sys_tmp736 = (w_sys_tmp737 + r_run_k_13);
	assign w_sys_tmp737 = 32'sh00000102;
	assign w_sys_tmp748 = (w_sys_tmp749 + r_run_k_13);
	assign w_sys_tmp749 = 32'sh00000121;
	assign w_sys_tmp760 = (w_sys_tmp761 + r_run_k_13);
	assign w_sys_tmp761 = 32'sh00000140;
	assign w_sys_tmp772 = (w_sys_tmp773 + r_run_k_13);
	assign w_sys_tmp773 = 32'sh0000015f;
	assign w_sys_tmp784 = (w_sys_tmp785 + r_run_k_13);
	assign w_sys_tmp785 = 32'sh0000017e;
	assign w_sys_tmp820 = (w_sys_tmp821 + r_run_k_13);
	assign w_sys_tmp821 = 32'sh0000019d;
	assign w_sys_tmp832 = (w_sys_tmp833 + r_run_k_13);
	assign w_sys_tmp833 = 32'sh000001bc;
	assign w_sys_tmp844 = (w_sys_tmp845 + r_run_k_13);
	assign w_sys_tmp845 = 32'sh000001db;
	assign w_sys_tmp856 = (w_sys_tmp857 + r_run_k_13);
	assign w_sys_tmp857 = 32'sh000001fa;
	assign w_sys_tmp868 = (w_sys_tmp869 + r_run_k_13);
	assign w_sys_tmp869 = 32'sh00000219;
	assign w_sys_tmp880 = (w_sys_tmp881 + r_run_k_13);
	assign w_sys_tmp881 = 32'sh00000238;
	assign w_sys_tmp892 = (w_sys_tmp893 + r_run_k_13);
	assign w_sys_tmp893 = 32'sh00000257;
	assign w_sys_tmp904 = (w_sys_tmp905 + r_run_k_13);
	assign w_sys_tmp905 = 32'sh00000276;
	assign w_sys_tmp916 = (w_sys_tmp917 + r_run_k_13);
	assign w_sys_tmp917 = 32'sh00000295;
	assign w_sys_tmp928 = (w_sys_tmp929 + r_run_k_13);
	assign w_sys_tmp929 = 32'sh000002b4;
	assign w_sys_tmp964 = (w_sys_tmp965 + r_run_k_13);
	assign w_sys_tmp965 = 32'sh000002d3;
	assign w_sys_tmp976 = (w_sys_tmp977 + r_run_k_13);
	assign w_sys_tmp977 = 32'sh000002f2;
	assign w_sys_tmp988 = (w_sys_tmp989 + r_run_k_13);
	assign w_sys_tmp989 = 32'sh00000311;
	assign w_sys_tmp1000 = (w_sys_tmp1001 + r_run_k_13);
	assign w_sys_tmp1001 = 32'sh00000330;
	assign w_sys_tmp1012 = (w_sys_tmp1013 + r_run_k_13);
	assign w_sys_tmp1013 = 32'sh0000034f;
	assign w_sys_tmp1024 = (w_sys_tmp1025 + r_run_k_13);
	assign w_sys_tmp1025 = 32'sh0000036e;
	assign w_sys_tmp1036 = (w_sys_tmp1037 + r_run_k_13);
	assign w_sys_tmp1037 = 32'sh0000038d;
	assign w_sys_tmp1048 = (w_sys_tmp1049 + r_run_k_13);
	assign w_sys_tmp1049 = 32'sh000003ac;
	assign w_sys_tmp1060 = (w_sys_tmp1061 + r_run_k_13);
	assign w_sys_tmp1061 = 32'sh000003cb;
	assign w_sys_tmp1071 = (r_run_k_13 + w_sys_intOne);
	assign w_sys_tmp1072 = 32'sh00000015;
	assign w_sys_tmp1073 = ( !w_sys_tmp1074 );
	assign w_sys_tmp1074 = (w_sys_tmp1075 < r_run_k_13);
	assign w_sys_tmp1075 = 32'sh0000001f;
	assign w_sys_tmp1078 = (w_sys_tmp1079 + r_run_k_13);
	assign w_sys_tmp1079 = 32'sh0000001f;
	assign w_sys_tmp1080 = w_fld_U_2_dataout_1;
	assign w_sys_tmp1086 = w_fld_V_3_dataout_1;
	assign w_sys_tmp1090 = (w_sys_tmp1091 + r_run_k_13);
	assign w_sys_tmp1091 = 32'sh0000003e;
	assign w_sys_tmp1102 = (w_sys_tmp1103 + r_run_k_13);
	assign w_sys_tmp1103 = 32'sh0000005d;
	assign w_sys_tmp1114 = (w_sys_tmp1115 + r_run_k_13);
	assign w_sys_tmp1115 = 32'sh0000007c;
	assign w_sys_tmp1126 = (w_sys_tmp1127 + r_run_k_13);
	assign w_sys_tmp1127 = 32'sh0000009b;
	assign w_sys_tmp1138 = (w_sys_tmp1139 + r_run_k_13);
	assign w_sys_tmp1139 = 32'sh000000ba;
	assign w_sys_tmp1150 = (w_sys_tmp1151 + r_run_k_13);
	assign w_sys_tmp1151 = 32'sh000000d9;
	assign w_sys_tmp1162 = (w_sys_tmp1163 + r_run_k_13);
	assign w_sys_tmp1163 = 32'sh000000f8;
	assign w_sys_tmp1174 = (w_sys_tmp1175 + r_run_k_13);
	assign w_sys_tmp1175 = 32'sh00000117;
	assign w_sys_tmp1186 = (w_sys_tmp1187 + r_run_k_13);
	assign w_sys_tmp1187 = 32'sh00000136;
	assign w_sys_tmp1198 = (w_sys_tmp1199 + r_run_k_13);
	assign w_sys_tmp1199 = 32'sh00000155;
	assign w_sys_tmp1210 = (w_sys_tmp1211 + r_run_k_13);
	assign w_sys_tmp1211 = 32'sh00000174;
	assign w_sys_tmp1246 = (w_sys_tmp1247 + r_run_k_13);
	assign w_sys_tmp1247 = 32'sh00000193;
	assign w_sys_tmp1258 = (w_sys_tmp1259 + r_run_k_13);
	assign w_sys_tmp1259 = 32'sh000001b2;
	assign w_sys_tmp1270 = (w_sys_tmp1271 + r_run_k_13);
	assign w_sys_tmp1271 = 32'sh000001d1;
	assign w_sys_tmp1282 = (w_sys_tmp1283 + r_run_k_13);
	assign w_sys_tmp1283 = 32'sh000001f0;
	assign w_sys_tmp1294 = (w_sys_tmp1295 + r_run_k_13);
	assign w_sys_tmp1295 = 32'sh0000020f;
	assign w_sys_tmp1306 = (w_sys_tmp1307 + r_run_k_13);
	assign w_sys_tmp1307 = 32'sh0000022e;
	assign w_sys_tmp1318 = (w_sys_tmp1319 + r_run_k_13);
	assign w_sys_tmp1319 = 32'sh0000024d;
	assign w_sys_tmp1330 = (w_sys_tmp1331 + r_run_k_13);
	assign w_sys_tmp1331 = 32'sh0000026c;
	assign w_sys_tmp1342 = (w_sys_tmp1343 + r_run_k_13);
	assign w_sys_tmp1343 = 32'sh0000028b;
	assign w_sys_tmp1366 = (w_sys_tmp1367 + r_run_k_13);
	assign w_sys_tmp1367 = 32'sh000002aa;
	assign w_sys_tmp1378 = (w_sys_tmp1379 + r_run_k_13);
	assign w_sys_tmp1379 = 32'sh000002c9;
	assign w_sys_tmp1390 = (w_sys_tmp1391 + r_run_k_13);
	assign w_sys_tmp1391 = 32'sh000002e8;
	assign w_sys_tmp1402 = (w_sys_tmp1403 + r_run_k_13);
	assign w_sys_tmp1403 = 32'sh00000307;
	assign w_sys_tmp1414 = (w_sys_tmp1415 + r_run_k_13);
	assign w_sys_tmp1415 = 32'sh00000326;
	assign w_sys_tmp1426 = (w_sys_tmp1427 + r_run_k_13);
	assign w_sys_tmp1427 = 32'sh00000345;
	assign w_sys_tmp1438 = (w_sys_tmp1439 + r_run_k_13);
	assign w_sys_tmp1439 = 32'sh00000364;
	assign w_sys_tmp1450 = (w_sys_tmp1451 + r_run_k_13);
	assign w_sys_tmp1451 = 32'sh00000383;
	assign w_sys_tmp1462 = (w_sys_tmp1463 + r_run_k_13);
	assign w_sys_tmp1463 = 32'sh000003a2;
	assign w_sys_tmp1473 = (r_run_k_13 + w_sys_intOne);
	assign w_sys_tmp1474 = ( !w_sys_tmp1475 );
	assign w_sys_tmp1475 = (r_run_nlast_28 < r_run_n_15);
	assign w_sys_tmp1476 = (r_run_n_15 + w_sys_intOne);
	assign w_sys_tmp1477 = ( !w_sys_tmp1478 );
	assign w_sys_tmp1478 = (r_run_my_17 < r_run_k_13);
	assign w_sys_tmp1481 = (w_sys_tmp1482 + r_run_k_13);
	assign w_sys_tmp1482 = 32'sh0000001f;
	assign w_sys_tmp1483 = 32'h0;
	assign w_sys_tmp1485 = (w_sys_tmp1486 + r_run_k_13);
	assign w_sys_tmp1486 = (r_run_mx_16 * w_sys_tmp1482);
	assign w_sys_tmp1488 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1489 = (w_sys_tmp1490 + r_run_k_13);
	assign w_sys_tmp1490 = (w_sys_tmp1491 * w_sys_tmp1482);
	assign w_sys_tmp1491 = (r_run_mx_16 - w_sys_intOne);
	assign w_sys_tmp1493 = (r_run_k_13 + w_sys_intOne);
	assign w_sys_tmp1494 = ( !w_sys_tmp1495 );
	assign w_sys_tmp1495 = (r_run_mx_16 < r_run_j_14);
	assign w_sys_tmp1498 = (w_sys_tmp1499 + w_sys_intOne);
	assign w_sys_tmp1499 = (r_run_j_14 * w_sys_tmp1500);
	assign w_sys_tmp1500 = 32'sh0000001f;
	assign w_sys_tmp1501 = 32'h0;
	assign w_sys_tmp1503 = (w_sys_tmp1504 + r_run_my_17);
	assign w_sys_tmp1504 = (r_run_copy0_j_32 * w_sys_tmp1500);
	assign w_sys_tmp1507 = (r_run_copy0_j_32 + w_sys_intOne);
	assign w_sys_tmp1508 = (r_run_j_14 + w_sys_intOne);
	assign w_sys_tmp1581 = (r_run_mx_16 / w_sys_tmp1582);
	assign w_sys_tmp1582 = 32'sh00000004;
	assign w_sys_tmp1583 = ( !w_sys_tmp1584 );
	assign w_sys_tmp1584 = (w_sys_tmp1585 < r_run_j_14);
	assign w_sys_tmp1585 = (r_run_mx_16 / w_sys_tmp1586);
	assign w_sys_tmp1586 = 32'sh00000002;
	assign w_sys_tmp1589 = (w_sys_tmp1590 + w_sys_intOne);
	assign w_sys_tmp1590 = (r_run_j_14 * w_sys_tmp1591);
	assign w_sys_tmp1591 = 32'sh0000001f;
	assign w_sys_tmp1592 = 32'h3f800000;
	assign w_sys_tmp1593 = (r_run_j_14 + w_sys_intOne);
	assign w_sys_tmp1630 = ( !w_sys_tmp1631 );
	assign w_sys_tmp1631 = (w_sys_tmp1632 < r_run_k_13);
	assign w_sys_tmp1632 = 32'sh0000000c;
	assign w_sys_tmp1635 = (w_sys_tmp1636 + r_run_k_13);
	assign w_sys_tmp1636 = 32'sh0000001f;
	assign w_sys_tmp1637 = w_fld_T_0_dataout_1;
	assign w_sys_tmp1641 = (w_sys_tmp1642 + r_run_k_13);
	assign w_sys_tmp1642 = 32'sh0000003e;
	assign w_sys_tmp1647 = (w_sys_tmp1648 + r_run_k_13);
	assign w_sys_tmp1648 = 32'sh0000005d;
	assign w_sys_tmp1653 = (w_sys_tmp1654 + r_run_k_13);
	assign w_sys_tmp1654 = 32'sh0000007c;
	assign w_sys_tmp1659 = (w_sys_tmp1660 + r_run_k_13);
	assign w_sys_tmp1660 = 32'sh0000009b;
	assign w_sys_tmp1665 = (w_sys_tmp1666 + r_run_k_13);
	assign w_sys_tmp1666 = 32'sh000000ba;
	assign w_sys_tmp1671 = (w_sys_tmp1672 + r_run_k_13);
	assign w_sys_tmp1672 = 32'sh000000d9;
	assign w_sys_tmp1677 = (w_sys_tmp1678 + r_run_k_13);
	assign w_sys_tmp1678 = 32'sh000000f8;
	assign w_sys_tmp1683 = (w_sys_tmp1684 + r_run_k_13);
	assign w_sys_tmp1684 = 32'sh00000117;
	assign w_sys_tmp1689 = (w_sys_tmp1690 + r_run_k_13);
	assign w_sys_tmp1690 = 32'sh00000136;
	assign w_sys_tmp1695 = (w_sys_tmp1696 + r_run_k_13);
	assign w_sys_tmp1696 = 32'sh00000155;
	assign w_sys_tmp1701 = (w_sys_tmp1702 + r_run_k_13);
	assign w_sys_tmp1702 = 32'sh00000174;
	assign w_sys_tmp1719 = (w_sys_tmp1720 + r_run_k_13);
	assign w_sys_tmp1720 = 32'sh00000193;
	assign w_sys_tmp1725 = (w_sys_tmp1726 + r_run_k_13);
	assign w_sys_tmp1726 = 32'sh000001b2;
	assign w_sys_tmp1731 = (w_sys_tmp1732 + r_run_k_13);
	assign w_sys_tmp1732 = 32'sh000001d1;
	assign w_sys_tmp1737 = (w_sys_tmp1738 + r_run_k_13);
	assign w_sys_tmp1738 = 32'sh000001f0;
	assign w_sys_tmp1743 = (w_sys_tmp1744 + r_run_k_13);
	assign w_sys_tmp1744 = 32'sh0000020f;
	assign w_sys_tmp1749 = (w_sys_tmp1750 + r_run_k_13);
	assign w_sys_tmp1750 = 32'sh0000022e;
	assign w_sys_tmp1755 = (w_sys_tmp1756 + r_run_k_13);
	assign w_sys_tmp1756 = 32'sh0000024d;
	assign w_sys_tmp1761 = (w_sys_tmp1762 + r_run_k_13);
	assign w_sys_tmp1762 = 32'sh0000026c;
	assign w_sys_tmp1767 = (w_sys_tmp1768 + r_run_k_13);
	assign w_sys_tmp1768 = 32'sh0000028b;
	assign w_sys_tmp1773 = (w_sys_tmp1774 + r_run_k_13);
	assign w_sys_tmp1774 = 32'sh000002aa;
	assign w_sys_tmp1791 = (w_sys_tmp1792 + r_run_k_13);
	assign w_sys_tmp1792 = 32'sh000002c9;
	assign w_sys_tmp1797 = (w_sys_tmp1798 + r_run_k_13);
	assign w_sys_tmp1798 = 32'sh000002e8;
	assign w_sys_tmp1803 = (w_sys_tmp1804 + r_run_k_13);
	assign w_sys_tmp1804 = 32'sh00000307;
	assign w_sys_tmp1809 = (w_sys_tmp1810 + r_run_k_13);
	assign w_sys_tmp1810 = 32'sh00000326;
	assign w_sys_tmp1815 = (w_sys_tmp1816 + r_run_k_13);
	assign w_sys_tmp1816 = 32'sh00000345;
	assign w_sys_tmp1821 = (w_sys_tmp1822 + r_run_k_13);
	assign w_sys_tmp1822 = 32'sh00000364;
	assign w_sys_tmp1827 = (w_sys_tmp1828 + r_run_k_13);
	assign w_sys_tmp1828 = 32'sh00000383;
	assign w_sys_tmp1833 = (w_sys_tmp1834 + r_run_k_13);
	assign w_sys_tmp1834 = 32'sh000003a2;
	assign w_sys_tmp1839 = (w_sys_tmp1840 + r_run_k_13);
	assign w_sys_tmp1840 = 32'sh000003c1;
	assign w_sys_tmp1845 = (w_sys_tmp1846 + r_run_k_13);
	assign w_sys_tmp1846 = 32'sh00000029;
	assign w_sys_tmp1851 = (w_sys_tmp1852 + r_run_k_13);
	assign w_sys_tmp1852 = 32'sh00000048;
	assign w_sys_tmp1857 = (w_sys_tmp1858 + r_run_k_13);
	assign w_sys_tmp1858 = 32'sh00000067;
	assign w_sys_tmp1863 = (w_sys_tmp1864 + r_run_k_13);
	assign w_sys_tmp1864 = 32'sh00000086;
	assign w_sys_tmp1869 = (w_sys_tmp1870 + r_run_k_13);
	assign w_sys_tmp1870 = 32'sh000000a5;
	assign w_sys_tmp1875 = (w_sys_tmp1876 + r_run_k_13);
	assign w_sys_tmp1876 = 32'sh000000c4;
	assign w_sys_tmp1881 = (w_sys_tmp1882 + r_run_k_13);
	assign w_sys_tmp1882 = 32'sh000000e3;
	assign w_sys_tmp1887 = (w_sys_tmp1888 + r_run_k_13);
	assign w_sys_tmp1888 = 32'sh00000102;
	assign w_sys_tmp1893 = (w_sys_tmp1894 + r_run_k_13);
	assign w_sys_tmp1894 = 32'sh00000121;
	assign w_sys_tmp1899 = (w_sys_tmp1900 + r_run_k_13);
	assign w_sys_tmp1900 = 32'sh00000140;
	assign w_sys_tmp1905 = (w_sys_tmp1906 + r_run_k_13);
	assign w_sys_tmp1906 = 32'sh0000015f;
	assign w_sys_tmp1911 = (w_sys_tmp1912 + r_run_k_13);
	assign w_sys_tmp1912 = 32'sh0000017e;
	assign w_sys_tmp1929 = (w_sys_tmp1930 + r_run_k_13);
	assign w_sys_tmp1930 = 32'sh0000019d;
	assign w_sys_tmp1935 = (w_sys_tmp1936 + r_run_k_13);
	assign w_sys_tmp1936 = 32'sh000001bc;
	assign w_sys_tmp1941 = (w_sys_tmp1942 + r_run_k_13);
	assign w_sys_tmp1942 = 32'sh000001db;
	assign w_sys_tmp1947 = (w_sys_tmp1948 + r_run_k_13);
	assign w_sys_tmp1948 = 32'sh000001fa;
	assign w_sys_tmp1953 = (w_sys_tmp1954 + r_run_k_13);
	assign w_sys_tmp1954 = 32'sh00000219;
	assign w_sys_tmp1959 = (w_sys_tmp1960 + r_run_k_13);
	assign w_sys_tmp1960 = 32'sh00000238;
	assign w_sys_tmp1965 = (w_sys_tmp1966 + r_run_k_13);
	assign w_sys_tmp1966 = 32'sh00000257;
	assign w_sys_tmp1971 = (w_sys_tmp1972 + r_run_k_13);
	assign w_sys_tmp1972 = 32'sh00000276;
	assign w_sys_tmp1977 = (w_sys_tmp1978 + r_run_k_13);
	assign w_sys_tmp1978 = 32'sh00000295;
	assign w_sys_tmp1983 = (w_sys_tmp1984 + r_run_k_13);
	assign w_sys_tmp1984 = 32'sh000002b4;
	assign w_sys_tmp2001 = (w_sys_tmp2002 + r_run_k_13);
	assign w_sys_tmp2002 = 32'sh000002d3;
	assign w_sys_tmp2007 = (w_sys_tmp2008 + r_run_k_13);
	assign w_sys_tmp2008 = 32'sh000002f2;
	assign w_sys_tmp2013 = (w_sys_tmp2014 + r_run_k_13);
	assign w_sys_tmp2014 = 32'sh00000311;
	assign w_sys_tmp2019 = (w_sys_tmp2020 + r_run_k_13);
	assign w_sys_tmp2020 = 32'sh00000330;
	assign w_sys_tmp2025 = (w_sys_tmp2026 + r_run_k_13);
	assign w_sys_tmp2026 = 32'sh0000034f;
	assign w_sys_tmp2031 = (w_sys_tmp2032 + r_run_k_13);
	assign w_sys_tmp2032 = 32'sh0000036e;
	assign w_sys_tmp2037 = (w_sys_tmp2038 + r_run_k_13);
	assign w_sys_tmp2038 = 32'sh0000038d;
	assign w_sys_tmp2043 = (w_sys_tmp2044 + r_run_k_13);
	assign w_sys_tmp2044 = 32'sh000003ac;
	assign w_sys_tmp2049 = (w_sys_tmp2050 + r_run_k_13);
	assign w_sys_tmp2050 = 32'sh000003cb;
	assign w_sys_tmp2054 = (r_run_k_13 + w_sys_intOne);
	assign w_sys_tmp2055 = 32'sh00000015;
	assign w_sys_tmp2056 = ( !w_sys_tmp2057 );
	assign w_sys_tmp2057 = (w_sys_tmp2058 < r_run_k_13);
	assign w_sys_tmp2058 = 32'sh0000001f;
	assign w_sys_tmp2061 = (w_sys_tmp2062 + r_run_k_13);
	assign w_sys_tmp2062 = 32'sh0000001f;
	assign w_sys_tmp2063 = w_fld_T_0_dataout_1;
	assign w_sys_tmp2067 = (w_sys_tmp2068 + r_run_k_13);
	assign w_sys_tmp2068 = 32'sh0000003e;
	assign w_sys_tmp2073 = (w_sys_tmp2074 + r_run_k_13);
	assign w_sys_tmp2074 = 32'sh0000005d;
	assign w_sys_tmp2079 = (w_sys_tmp2080 + r_run_k_13);
	assign w_sys_tmp2080 = 32'sh0000007c;
	assign w_sys_tmp2085 = (w_sys_tmp2086 + r_run_k_13);
	assign w_sys_tmp2086 = 32'sh0000009b;
	assign w_sys_tmp2091 = (w_sys_tmp2092 + r_run_k_13);
	assign w_sys_tmp2092 = 32'sh000000ba;
	assign w_sys_tmp2097 = (w_sys_tmp2098 + r_run_k_13);
	assign w_sys_tmp2098 = 32'sh000000d9;
	assign w_sys_tmp2103 = (w_sys_tmp2104 + r_run_k_13);
	assign w_sys_tmp2104 = 32'sh000000f8;
	assign w_sys_tmp2109 = (w_sys_tmp2110 + r_run_k_13);
	assign w_sys_tmp2110 = 32'sh00000117;
	assign w_sys_tmp2115 = (w_sys_tmp2116 + r_run_k_13);
	assign w_sys_tmp2116 = 32'sh00000136;
	assign w_sys_tmp2121 = (w_sys_tmp2122 + r_run_k_13);
	assign w_sys_tmp2122 = 32'sh00000155;
	assign w_sys_tmp2127 = (w_sys_tmp2128 + r_run_k_13);
	assign w_sys_tmp2128 = 32'sh00000174;
	assign w_sys_tmp2145 = (w_sys_tmp2146 + r_run_k_13);
	assign w_sys_tmp2146 = 32'sh00000193;
	assign w_sys_tmp2151 = (w_sys_tmp2152 + r_run_k_13);
	assign w_sys_tmp2152 = 32'sh000001b2;
	assign w_sys_tmp2157 = (w_sys_tmp2158 + r_run_k_13);
	assign w_sys_tmp2158 = 32'sh000001d1;
	assign w_sys_tmp2163 = (w_sys_tmp2164 + r_run_k_13);
	assign w_sys_tmp2164 = 32'sh000001f0;
	assign w_sys_tmp2169 = (w_sys_tmp2170 + r_run_k_13);
	assign w_sys_tmp2170 = 32'sh0000020f;
	assign w_sys_tmp2175 = (w_sys_tmp2176 + r_run_k_13);
	assign w_sys_tmp2176 = 32'sh0000022e;
	assign w_sys_tmp2181 = (w_sys_tmp2182 + r_run_k_13);
	assign w_sys_tmp2182 = 32'sh0000024d;
	assign w_sys_tmp2187 = (w_sys_tmp2188 + r_run_k_13);
	assign w_sys_tmp2188 = 32'sh0000026c;
	assign w_sys_tmp2193 = (w_sys_tmp2194 + r_run_k_13);
	assign w_sys_tmp2194 = 32'sh0000028b;
	assign w_sys_tmp2199 = (w_sys_tmp2200 + r_run_k_13);
	assign w_sys_tmp2200 = 32'sh000002aa;
	assign w_sys_tmp2217 = (w_sys_tmp2218 + r_run_k_13);
	assign w_sys_tmp2218 = 32'sh000002c9;
	assign w_sys_tmp2223 = (w_sys_tmp2224 + r_run_k_13);
	assign w_sys_tmp2224 = 32'sh000002e8;
	assign w_sys_tmp2229 = (w_sys_tmp2230 + r_run_k_13);
	assign w_sys_tmp2230 = 32'sh00000307;
	assign w_sys_tmp2235 = (w_sys_tmp2236 + r_run_k_13);
	assign w_sys_tmp2236 = 32'sh00000345;
	assign w_sys_tmp2241 = (w_sys_tmp2242 + r_run_k_13);
	assign w_sys_tmp2242 = 32'sh00000364;
	assign w_sys_tmp2247 = (w_sys_tmp2248 + r_run_k_13);
	assign w_sys_tmp2248 = 32'sh00000383;
	assign w_sys_tmp2253 = (w_sys_tmp2254 + r_run_k_13);
	assign w_sys_tmp2254 = 32'sh000003a2;
	assign w_sys_tmp2259 = (w_sys_tmp2260 + r_run_k_13);
	assign w_sys_tmp2260 = 32'sh000003c1;
	assign w_sys_tmp2264 = (r_run_k_13 + w_sys_intOne);
	assign w_sys_tmp2265 = 32'sh00000002;
	assign w_sys_tmp2266 = ( !w_sys_tmp2267 );
	assign w_sys_tmp2267 = (w_sys_tmp2268 < r_run_k_13);
	assign w_sys_tmp2268 = 32'sh0000000b;
	assign w_sys_tmp2271 = (w_sys_tmp2272 + r_run_k_13);
	assign w_sys_tmp2272 = 32'sh0000003e;
	assign w_sys_tmp2273 = w_sub00_result_dataout;
	assign w_sys_tmp2277 = (w_sys_tmp2278 + r_run_k_13);
	assign w_sys_tmp2278 = 32'sh0000005d;
	assign w_sys_tmp2283 = (w_sys_tmp2284 + r_run_k_13);
	assign w_sys_tmp2284 = 32'sh0000007c;
	assign w_sys_tmp2289 = (w_sys_tmp2290 + r_run_k_13);
	assign w_sys_tmp2290 = 32'sh0000009b;
	assign w_sys_tmp2295 = (w_sys_tmp2296 + r_run_k_13);
	assign w_sys_tmp2296 = 32'sh000000ba;
	assign w_sys_tmp2301 = (w_sys_tmp2302 + r_run_k_13);
	assign w_sys_tmp2302 = 32'sh000000d9;
	assign w_sys_tmp2307 = (w_sys_tmp2308 + r_run_k_13);
	assign w_sys_tmp2308 = 32'sh000000f8;
	assign w_sys_tmp2313 = (w_sys_tmp2314 + r_run_k_13);
	assign w_sys_tmp2314 = 32'sh00000117;
	assign w_sys_tmp2319 = (w_sys_tmp2320 + r_run_k_13);
	assign w_sys_tmp2320 = 32'sh00000136;
	assign w_sys_tmp2325 = (w_sys_tmp2326 + r_run_k_13);
	assign w_sys_tmp2326 = 32'sh00000155;
	assign w_sys_tmp2331 = (w_sys_tmp2332 + r_run_k_13);
	assign w_sys_tmp2332 = 32'sh00000174;
	assign w_sys_tmp2336 = (w_sys_tmp2337 + r_run_k_13);
	assign w_sys_tmp2337 = 32'sh00000193;
	assign w_sys_tmp2341 = (w_sys_tmp2342 + r_run_k_13);
	assign w_sys_tmp2342 = 32'sh000001b2;
	assign w_sys_tmp2346 = (w_sys_tmp2347 + r_run_k_13);
	assign w_sys_tmp2347 = 32'sh000001d1;
	assign w_sys_tmp2351 = (w_sys_tmp2352 + r_run_k_13);
	assign w_sys_tmp2352 = 32'sh000001f0;
	assign w_sys_tmp2356 = (w_sys_tmp2357 + r_run_k_13);
	assign w_sys_tmp2357 = 32'sh0000020f;
	assign w_sys_tmp2361 = (w_sys_tmp2362 + r_run_k_13);
	assign w_sys_tmp2362 = 32'sh0000022e;
	assign w_sys_tmp2366 = (w_sys_tmp2367 + r_run_k_13);
	assign w_sys_tmp2367 = 32'sh0000024d;
	assign w_sys_tmp2371 = (w_sys_tmp2372 + r_run_k_13);
	assign w_sys_tmp2372 = 32'sh0000026c;
	assign w_sys_tmp2376 = (w_sys_tmp2377 + r_run_k_13);
	assign w_sys_tmp2377 = 32'sh0000028b;
	assign w_sys_tmp2381 = (w_sys_tmp2382 + r_run_k_13);
	assign w_sys_tmp2382 = 32'sh000002aa;
	assign w_sys_tmp2386 = (w_sys_tmp2387 + r_run_k_13);
	assign w_sys_tmp2387 = 32'sh000002c9;
	assign w_sys_tmp2391 = (w_sys_tmp2392 + r_run_k_13);
	assign w_sys_tmp2392 = 32'sh000002e8;
	assign w_sys_tmp2396 = (w_sys_tmp2397 + r_run_k_13);
	assign w_sys_tmp2397 = 32'sh00000307;
	assign w_sys_tmp2401 = (w_sys_tmp2402 + r_run_k_13);
	assign w_sys_tmp2402 = 32'sh00000326;
	assign w_sys_tmp2406 = (w_sys_tmp2407 + r_run_k_13);
	assign w_sys_tmp2407 = 32'sh00000345;
	assign w_sys_tmp2411 = (w_sys_tmp2412 + r_run_k_13);
	assign w_sys_tmp2412 = 32'sh00000364;
	assign w_sys_tmp2416 = (w_sys_tmp2417 + r_run_k_13);
	assign w_sys_tmp2417 = 32'sh00000383;
	assign w_sys_tmp2421 = (w_sys_tmp2422 + r_run_k_13);
	assign w_sys_tmp2422 = 32'sh000003a2;
	assign w_sys_tmp2426 = (w_sys_tmp2427 + r_run_k_13);
	assign w_sys_tmp2427 = 32'sh00000048;
	assign w_sys_tmp2431 = (w_sys_tmp2432 + r_run_k_13);
	assign w_sys_tmp2432 = 32'sh00000067;
	assign w_sys_tmp2436 = (w_sys_tmp2437 + r_run_k_13);
	assign w_sys_tmp2437 = 32'sh00000086;
	assign w_sys_tmp2441 = (w_sys_tmp2442 + r_run_k_13);
	assign w_sys_tmp2442 = 32'sh000000a5;
	assign w_sys_tmp2446 = (w_sys_tmp2447 + r_run_k_13);
	assign w_sys_tmp2447 = 32'sh000000c4;
	assign w_sys_tmp2451 = (w_sys_tmp2452 + r_run_k_13);
	assign w_sys_tmp2452 = 32'sh000000e3;
	assign w_sys_tmp2456 = (w_sys_tmp2457 + r_run_k_13);
	assign w_sys_tmp2457 = 32'sh00000102;
	assign w_sys_tmp2461 = (w_sys_tmp2462 + r_run_k_13);
	assign w_sys_tmp2462 = 32'sh00000121;
	assign w_sys_tmp2466 = (w_sys_tmp2467 + r_run_k_13);
	assign w_sys_tmp2467 = 32'sh00000140;
	assign w_sys_tmp2471 = (w_sys_tmp2472 + r_run_k_13);
	assign w_sys_tmp2472 = 32'sh0000015f;
	assign w_sys_tmp2476 = (w_sys_tmp2477 + r_run_k_13);
	assign w_sys_tmp2477 = 32'sh0000017e;
	assign w_sys_tmp2481 = (w_sys_tmp2482 + r_run_k_13);
	assign w_sys_tmp2482 = 32'sh0000019d;
	assign w_sys_tmp2486 = (w_sys_tmp2487 + r_run_k_13);
	assign w_sys_tmp2487 = 32'sh000001bc;
	assign w_sys_tmp2491 = (w_sys_tmp2492 + r_run_k_13);
	assign w_sys_tmp2492 = 32'sh000001db;
	assign w_sys_tmp2496 = (w_sys_tmp2497 + r_run_k_13);
	assign w_sys_tmp2497 = 32'sh000001fa;
	assign w_sys_tmp2501 = (w_sys_tmp2502 + r_run_k_13);
	assign w_sys_tmp2502 = 32'sh00000219;
	assign w_sys_tmp2506 = (w_sys_tmp2507 + r_run_k_13);
	assign w_sys_tmp2507 = 32'sh00000238;
	assign w_sys_tmp2511 = (w_sys_tmp2512 + r_run_k_13);
	assign w_sys_tmp2512 = 32'sh00000257;
	assign w_sys_tmp2516 = (w_sys_tmp2517 + r_run_k_13);
	assign w_sys_tmp2517 = 32'sh00000276;
	assign w_sys_tmp2521 = (w_sys_tmp2522 + r_run_k_13);
	assign w_sys_tmp2522 = 32'sh00000295;
	assign w_sys_tmp2526 = (w_sys_tmp2527 + r_run_k_13);
	assign w_sys_tmp2527 = 32'sh000002b4;
	assign w_sys_tmp2531 = (w_sys_tmp2532 + r_run_k_13);
	assign w_sys_tmp2532 = 32'sh000002d3;
	assign w_sys_tmp2536 = (w_sys_tmp2537 + r_run_k_13);
	assign w_sys_tmp2537 = 32'sh000002f2;
	assign w_sys_tmp2541 = (w_sys_tmp2542 + r_run_k_13);
	assign w_sys_tmp2542 = 32'sh00000311;
	assign w_sys_tmp2546 = (w_sys_tmp2547 + r_run_k_13);
	assign w_sys_tmp2547 = 32'sh00000330;
	assign w_sys_tmp2551 = (w_sys_tmp2552 + r_run_k_13);
	assign w_sys_tmp2552 = 32'sh0000034f;
	assign w_sys_tmp2556 = (w_sys_tmp2557 + r_run_k_13);
	assign w_sys_tmp2557 = 32'sh0000036e;
	assign w_sys_tmp2561 = (w_sys_tmp2562 + r_run_k_13);
	assign w_sys_tmp2562 = 32'sh0000038d;
	assign w_sys_tmp2566 = (w_sys_tmp2567 + r_run_k_13);
	assign w_sys_tmp2567 = 32'sh000003ac;
	assign w_sys_tmp2570 = (r_run_k_13 + w_sys_intOne);
	assign w_sys_tmp2571 = 32'sh00000016;
	assign w_sys_tmp2572 = ( !w_sys_tmp2573 );
	assign w_sys_tmp2573 = (w_sys_tmp2574 < r_run_k_13);
	assign w_sys_tmp2574 = 32'sh0000001e;
	assign w_sys_tmp2577 = (w_sys_tmp2578 + r_run_k_13);
	assign w_sys_tmp2578 = 32'sh0000003e;
	assign w_sys_tmp2579 = w_sub06_result_dataout;
	assign w_sys_tmp2583 = (w_sys_tmp2584 + r_run_k_13);
	assign w_sys_tmp2584 = 32'sh0000005d;
	assign w_sys_tmp2589 = (w_sys_tmp2590 + r_run_k_13);
	assign w_sys_tmp2590 = 32'sh0000007c;
	assign w_sys_tmp2595 = (w_sys_tmp2596 + r_run_k_13);
	assign w_sys_tmp2596 = 32'sh0000009b;
	assign w_sys_tmp2601 = (w_sys_tmp2602 + r_run_k_13);
	assign w_sys_tmp2602 = 32'sh000000ba;
	assign w_sys_tmp2607 = (w_sys_tmp2608 + r_run_k_13);
	assign w_sys_tmp2608 = 32'sh000000d9;
	assign w_sys_tmp2613 = (w_sys_tmp2614 + r_run_k_13);
	assign w_sys_tmp2614 = 32'sh000000f8;
	assign w_sys_tmp2619 = (w_sys_tmp2620 + r_run_k_13);
	assign w_sys_tmp2620 = 32'sh00000117;
	assign w_sys_tmp2625 = (w_sys_tmp2626 + r_run_k_13);
	assign w_sys_tmp2626 = 32'sh00000136;
	assign w_sys_tmp2631 = (w_sys_tmp2632 + r_run_k_13);
	assign w_sys_tmp2632 = 32'sh00000155;
	assign w_sys_tmp2637 = (w_sys_tmp2638 + r_run_k_13);
	assign w_sys_tmp2638 = 32'sh00000174;
	assign w_sys_tmp2642 = (w_sys_tmp2643 + r_run_k_13);
	assign w_sys_tmp2643 = 32'sh00000193;
	assign w_sys_tmp2647 = (w_sys_tmp2648 + r_run_k_13);
	assign w_sys_tmp2648 = 32'sh000001b2;
	assign w_sys_tmp2652 = (w_sys_tmp2653 + r_run_k_13);
	assign w_sys_tmp2653 = 32'sh000001d1;
	assign w_sys_tmp2657 = (w_sys_tmp2658 + r_run_k_13);
	assign w_sys_tmp2658 = 32'sh000001f0;
	assign w_sys_tmp2662 = (w_sys_tmp2663 + r_run_k_13);
	assign w_sys_tmp2663 = 32'sh0000020f;
	assign w_sys_tmp2667 = (w_sys_tmp2668 + r_run_k_13);
	assign w_sys_tmp2668 = 32'sh0000022e;
	assign w_sys_tmp2672 = (w_sys_tmp2673 + r_run_k_13);
	assign w_sys_tmp2673 = 32'sh0000024d;
	assign w_sys_tmp2677 = (w_sys_tmp2678 + r_run_k_13);
	assign w_sys_tmp2678 = 32'sh0000026c;
	assign w_sys_tmp2682 = (w_sys_tmp2683 + r_run_k_13);
	assign w_sys_tmp2683 = 32'sh0000028b;
	assign w_sys_tmp2687 = (w_sys_tmp2688 + r_run_k_13);
	assign w_sys_tmp2688 = 32'sh000002aa;
	assign w_sys_tmp2692 = (w_sys_tmp2693 + r_run_k_13);
	assign w_sys_tmp2693 = 32'sh000002c9;
	assign w_sys_tmp2697 = (w_sys_tmp2698 + r_run_k_13);
	assign w_sys_tmp2698 = 32'sh000002e8;
	assign w_sys_tmp2702 = (w_sys_tmp2703 + r_run_k_13);
	assign w_sys_tmp2703 = 32'sh00000307;
	assign w_sys_tmp2707 = (w_sys_tmp2708 + r_run_k_13);
	assign w_sys_tmp2708 = 32'sh00000326;
	assign w_sys_tmp2712 = (w_sys_tmp2713 + r_run_k_13);
	assign w_sys_tmp2713 = 32'sh00000345;
	assign w_sys_tmp2717 = (w_sys_tmp2718 + r_run_k_13);
	assign w_sys_tmp2718 = 32'sh00000364;
	assign w_sys_tmp2722 = (w_sys_tmp2723 + r_run_k_13);
	assign w_sys_tmp2723 = 32'sh00000383;
	assign w_sys_tmp2727 = (w_sys_tmp2728 + r_run_k_13);
	assign w_sys_tmp2728 = 32'sh000003a2;
	assign w_sys_tmp2731 = (r_run_k_13 + w_sys_intOne);


	sub08
		sub08_inst(
			.i_fld_T_0_addr_0 (w_sub08_T_addr),
			.i_fld_T_0_datain_0 (w_sub08_T_datain),
			.o_fld_T_0_dataout_0 (w_sub08_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub08_T_r_w),
			.i_fld_U_2_addr_0 (w_sub08_U_addr),
			.i_fld_U_2_datain_0 (w_sub08_U_datain),
			.o_fld_U_2_dataout_0 (w_sub08_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub08_U_r_w),
			.i_fld_V_1_addr_0 (w_sub08_V_addr),
			.i_fld_V_1_datain_0 (w_sub08_V_datain),
			.o_fld_V_1_dataout_0 (w_sub08_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub08_V_r_w),
			.i_fld_result_3_addr_0 (w_sub08_result_addr),
			.i_fld_result_3_datain_0 (w_sub08_result_datain),
			.o_fld_result_3_dataout_0 (w_sub08_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub08_result_r_w),
			.o_run_busy (w_sub08_run_busy),
			.i_run_req (r_sub08_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub03
		sub03_inst(
			.i_fld_T_0_addr_0 (w_sub03_T_addr),
			.i_fld_T_0_datain_0 (w_sub03_T_datain),
			.o_fld_T_0_dataout_0 (w_sub03_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub03_T_r_w),
			.i_fld_U_2_addr_0 (w_sub03_U_addr),
			.i_fld_U_2_datain_0 (w_sub03_U_datain),
			.o_fld_U_2_dataout_0 (w_sub03_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub03_U_r_w),
			.i_fld_V_1_addr_0 (w_sub03_V_addr),
			.i_fld_V_1_datain_0 (w_sub03_V_datain),
			.o_fld_V_1_dataout_0 (w_sub03_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub03_V_r_w),
			.i_fld_result_3_addr_0 (w_sub03_result_addr),
			.i_fld_result_3_datain_0 (w_sub03_result_datain),
			.o_fld_result_3_dataout_0 (w_sub03_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub03_result_r_w),
			.o_run_busy (w_sub03_run_busy),
			.i_run_req (r_sub03_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub02
		sub02_inst(
			.i_fld_T_0_addr_0 (w_sub02_T_addr),
			.i_fld_T_0_datain_0 (w_sub02_T_datain),
			.o_fld_T_0_dataout_0 (w_sub02_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub02_T_r_w),
			.i_fld_U_2_addr_0 (w_sub02_U_addr),
			.i_fld_U_2_datain_0 (w_sub02_U_datain),
			.o_fld_U_2_dataout_0 (w_sub02_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub02_U_r_w),
			.i_fld_V_1_addr_0 (w_sub02_V_addr),
			.i_fld_V_1_datain_0 (w_sub02_V_datain),
			.o_fld_V_1_dataout_0 (w_sub02_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub02_V_r_w),
			.i_fld_result_3_addr_0 (w_sub02_result_addr),
			.i_fld_result_3_datain_0 (w_sub02_result_datain),
			.o_fld_result_3_dataout_0 (w_sub02_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub02_result_r_w),
			.o_run_busy (w_sub02_run_busy),
			.i_run_req (r_sub02_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub01
		sub01_inst(
			.i_fld_T_0_addr_0 (w_sub01_T_addr),
			.i_fld_T_0_datain_0 (w_sub01_T_datain),
			.o_fld_T_0_dataout_0 (w_sub01_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub01_T_r_w),
			.i_fld_U_2_addr_0 (w_sub01_U_addr),
			.i_fld_U_2_datain_0 (w_sub01_U_datain),
			.o_fld_U_2_dataout_0 (w_sub01_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub01_U_r_w),
			.i_fld_V_1_addr_0 (w_sub01_V_addr),
			.i_fld_V_1_datain_0 (w_sub01_V_datain),
			.o_fld_V_1_dataout_0 (w_sub01_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub01_V_r_w),
			.i_fld_result_3_addr_0 (w_sub01_result_addr),
			.i_fld_result_3_datain_0 (w_sub01_result_datain),
			.o_fld_result_3_dataout_0 (w_sub01_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub01_result_r_w),
			.o_run_busy (w_sub01_run_busy),
			.i_run_req (r_sub01_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub00
		sub00_inst(
			.i_fld_T_0_addr_0 (w_sub00_T_addr),
			.i_fld_T_0_datain_0 (w_sub00_T_datain),
			.o_fld_T_0_dataout_0 (w_sub00_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub00_T_r_w),
			.i_fld_U_2_addr_0 (w_sub00_U_addr),
			.i_fld_U_2_datain_0 (w_sub00_U_datain),
			.o_fld_U_2_dataout_0 (w_sub00_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub00_U_r_w),
			.i_fld_V_1_addr_0 (w_sub00_V_addr),
			.i_fld_V_1_datain_0 (w_sub00_V_datain),
			.o_fld_V_1_dataout_0 (w_sub00_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub00_V_r_w),
			.i_fld_result_3_addr_0 (w_sub00_result_addr),
			.i_fld_result_3_datain_0 (w_sub00_result_datain),
			.o_fld_result_3_dataout_0 (w_sub00_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub00_result_r_w),
			.o_run_busy (w_sub00_run_busy),
			.i_run_req (r_sub00_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub07
		sub07_inst(
			.i_fld_T_0_addr_0 (w_sub07_T_addr),
			.i_fld_T_0_datain_0 (w_sub07_T_datain),
			.o_fld_T_0_dataout_0 (w_sub07_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub07_T_r_w),
			.i_fld_U_2_addr_0 (w_sub07_U_addr),
			.i_fld_U_2_datain_0 (w_sub07_U_datain),
			.o_fld_U_2_dataout_0 (w_sub07_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub07_U_r_w),
			.i_fld_V_1_addr_0 (w_sub07_V_addr),
			.i_fld_V_1_datain_0 (w_sub07_V_datain),
			.o_fld_V_1_dataout_0 (w_sub07_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub07_V_r_w),
			.i_fld_result_3_addr_0 (w_sub07_result_addr),
			.i_fld_result_3_datain_0 (w_sub07_result_datain),
			.o_fld_result_3_dataout_0 (w_sub07_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub07_result_r_w),
			.o_run_busy (w_sub07_run_busy),
			.i_run_req (r_sub07_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub06
		sub06_inst(
			.i_fld_T_0_addr_0 (w_sub06_T_addr),
			.i_fld_T_0_datain_0 (w_sub06_T_datain),
			.o_fld_T_0_dataout_0 (w_sub06_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub06_T_r_w),
			.i_fld_U_2_addr_0 (w_sub06_U_addr),
			.i_fld_U_2_datain_0 (w_sub06_U_datain),
			.o_fld_U_2_dataout_0 (w_sub06_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub06_U_r_w),
			.i_fld_V_1_addr_0 (w_sub06_V_addr),
			.i_fld_V_1_datain_0 (w_sub06_V_datain),
			.o_fld_V_1_dataout_0 (w_sub06_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub06_V_r_w),
			.i_fld_result_3_addr_0 (w_sub06_result_addr),
			.i_fld_result_3_datain_0 (w_sub06_result_datain),
			.o_fld_result_3_dataout_0 (w_sub06_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub06_result_r_w),
			.o_run_busy (w_sub06_run_busy),
			.i_run_req (r_sub06_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub05
		sub05_inst(
			.i_fld_T_0_addr_0 (w_sub05_T_addr),
			.i_fld_T_0_datain_0 (w_sub05_T_datain),
			.o_fld_T_0_dataout_0 (w_sub05_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub05_T_r_w),
			.i_fld_U_2_addr_0 (w_sub05_U_addr),
			.i_fld_U_2_datain_0 (w_sub05_U_datain),
			.o_fld_U_2_dataout_0 (w_sub05_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub05_U_r_w),
			.i_fld_V_1_addr_0 (w_sub05_V_addr),
			.i_fld_V_1_datain_0 (w_sub05_V_datain),
			.o_fld_V_1_dataout_0 (w_sub05_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub05_V_r_w),
			.i_fld_result_3_addr_0 (w_sub05_result_addr),
			.i_fld_result_3_datain_0 (w_sub05_result_datain),
			.o_fld_result_3_dataout_0 (w_sub05_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub05_result_r_w),
			.o_run_busy (w_sub05_run_busy),
			.i_run_req (r_sub05_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	sub04
		sub04_inst(
			.i_fld_T_0_addr_0 (w_sub04_T_addr),
			.i_fld_T_0_datain_0 (w_sub04_T_datain),
			.o_fld_T_0_dataout_0 (w_sub04_T_dataout),
			.i_fld_T_0_r_w_0 (w_sub04_T_r_w),
			.i_fld_U_2_addr_0 (w_sub04_U_addr),
			.i_fld_U_2_datain_0 (w_sub04_U_datain),
			.o_fld_U_2_dataout_0 (w_sub04_U_dataout),
			.i_fld_U_2_r_w_0 (w_sub04_U_r_w),
			.i_fld_V_1_addr_0 (w_sub04_V_addr),
			.i_fld_V_1_datain_0 (w_sub04_V_datain),
			.o_fld_V_1_dataout_0 (w_sub04_V_dataout),
			.i_fld_V_1_r_w_0 (w_sub04_V_r_w),
			.i_fld_result_3_addr_0 (w_sub04_result_addr),
			.i_fld_result_3_datain_0 (w_sub04_result_datain),
			.o_fld_result_3_dataout_0 (w_sub04_result_dataout),
			.i_fld_result_3_r_w_0 (w_sub04_result_r_w),
			.o_run_busy (w_sub04_run_busy),
			.i_run_req (r_sub04_run_req),
			.ce (ce),
			.reset_n (reset_n),
			.clock (clock)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_T_0(
			.clk (clock),
			.ce_0 (w_fld_T_0_ce_0),
			.addr_0 (w_fld_T_0_addr_0),
			.datain_0 (w_fld_T_0_datain_0),
			.dataout_0 (w_fld_T_0_dataout_0),
			.r_w_0 (w_fld_T_0_r_w_0),
			.ce_1 (w_fld_T_0_ce_1),
			.addr_1 (r_fld_T_0_addr_1),
			.datain_1 (r_fld_T_0_datain_1),
			.dataout_1 (w_fld_T_0_dataout_1),
			.r_w_1 (r_fld_T_0_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_TT_1(
			.clk (clock),
			.ce_0 (w_fld_TT_1_ce_0),
			.addr_0 (w_fld_TT_1_addr_0),
			.datain_0 (w_fld_TT_1_datain_0),
			.dataout_0 (w_fld_TT_1_dataout_0),
			.r_w_0 (w_fld_TT_1_r_w_0),
			.ce_1 (w_fld_TT_1_ce_1),
			.addr_1 (r_fld_TT_1_addr_1),
			.datain_1 (r_fld_TT_1_datain_1),
			.dataout_1 (w_fld_TT_1_dataout_1),
			.r_w_1 (r_fld_TT_1_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_U_2(
			.clk (clock),
			.ce_0 (w_fld_U_2_ce_0),
			.addr_0 (w_fld_U_2_addr_0),
			.datain_0 (w_fld_U_2_datain_0),
			.dataout_0 (w_fld_U_2_dataout_0),
			.r_w_0 (w_fld_U_2_r_w_0),
			.ce_1 (w_fld_U_2_ce_1),
			.addr_1 (r_fld_U_2_addr_1),
			.datain_1 (r_fld_U_2_datain_1),
			.dataout_1 (w_fld_U_2_dataout_1),
			.r_w_1 (r_fld_U_2_r_w_1)
		);

	DualPortRAM #(.DWIDTH(32), .AWIDTH(9), .WORDS(484) )
		dpram_V_3(
			.clk (clock),
			.ce_0 (w_fld_V_3_ce_0),
			.addr_0 (w_fld_V_3_addr_0),
			.datain_0 (w_fld_V_3_datain_0),
			.dataout_0 (w_fld_V_3_dataout_0),
			.r_w_0 (w_fld_V_3_r_w_0),
			.ce_1 (w_fld_V_3_ce_1),
			.addr_1 (r_fld_V_3_addr_1),
			.datain_1 (r_fld_V_3_datain_1),
			.dataout_1 (w_fld_V_3_dataout_1),
			.r_w_1 (r_fld_V_3_r_w_1)
		);

	AddFloat
		AddFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_AddFloat_portA_0),
			.b (r_ip_AddFloat_portB_0),
			.result (w_ip_AddFloat_result_0)
		);

	MultFloat
		MultFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_MultFloat_multiplicand_0),
			.b (r_ip_MultFloat_multiplier_0),
			.result (w_ip_MultFloat_product_0)
		);

	FixedToFloat
		FixedToFloat_inst_0(
			.clk (clock),
			.ce (w_sys_ce),
			.a (r_ip_FixedToFloat_fixed_0),
			.result (w_ip_FixedToFloat_floating_0)
		);

	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14)) begin
										r_ip_AddFloat_portA_0 <= w_sys_tmp39;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp129[31], w_sys_tmp129[30:0] };

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp129[31], w_sys_tmp129[30:0] };

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_ip_AddFloat_portB_0 <= { ~w_sys_tmp38[31], w_sys_tmp38[30:0] };

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h18)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19) || (r_sys_run_step==7'h1a)) begin
										r_ip_MultFloat_multiplicand_0 <= r_sys_tmp4_float;

									end
									else
									if((7'h7<=r_sys_run_step && r_sys_run_step<=7'hb) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'hf)) begin
										r_ip_MultFloat_multiplicand_0 <= r_run_dy_20;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp19;

									end
									else
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h16)) begin
										r_ip_MultFloat_multiplicand_0 <= w_sys_tmp37;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'he) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14) || (r_sys_run_step==7'h16)) begin
										r_ip_MultFloat_multiplier_0 <= r_run_YY_25;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp38;

									end
									else
									if((r_sys_run_step==7'h15) || (r_sys_run_step==7'h18) || (r_sys_run_step==7'h1b)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp2_float;

									end
									else
									if((7'h7<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_ip_MultFloat_multiplier_0 <= w_sys_tmp20;

									end
									else
									if((r_sys_run_step==7'hd) || (r_sys_run_step==7'hf)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h13) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h1a)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_ip_MultFloat_multiplier_0 <= r_sys_tmp1_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_ip_FixedToFloat_fixed_0 <= w_sys_tmp21;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_processing_methodID <= 2'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_processing_methodID <= ((i_run_req) ? 2'h1 : r_sys_processing_methodID);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h4d: begin
							r_sys_processing_methodID <= r_sys_run_caller;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_caller <= 2'h0;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_req <= w_sys_boolFalse;

		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_phase <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_phase <= 7'h2;
						end

						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h4;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp13) ? 7'h9 : 7'hf);

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h5;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp16) ? 7'hd : 7'h6);

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h20)) begin
										r_sys_run_phase <= 7'ha;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp227) ? 7'h13 : 7'h15);

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_phase <= 7'h10;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1073) ? 7'h19 : 7'h1b);

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sys_run_phase <= 7'h16;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1474) ? 7'h20 : 7'h4d);

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h1c;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1477) ? 7'h24 : 7'h26);

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_run_phase <= 7'h21;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1494) ? 7'h2a : 7'h2c);

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_phase <= 7'h27;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1583) ? 7'h30 : 7'h32);

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_phase <= 7'h2d;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp1630) ? 7'h36 : 7'h38);

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_phase <= 7'h33;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2056) ? 7'h3c : 7'h3d);

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h23)) begin
										r_sys_run_phase <= 7'h39;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 7'h3f;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_phase <= 7'h41;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h42;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2266) ? 7'h45 : 7'h47);

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3b)) begin
										r_sys_run_phase <= 7'h42;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= 7'h48;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_phase <= ((w_sys_tmp2572) ? 7'h4b : 7'h1d);

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_sys_run_phase <= 7'h48;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sys_run_phase <= 7'h0;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_stage <= 4'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h20)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h23)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= w_sys_run_stage_p1;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3b)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_sys_run_stage <= 4'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_step <= 7'h0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h5: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'ha: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h20)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1f)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h10: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h46)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h16: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h21)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h21: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h1) || (r_sys_run_step==7'h2)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h27: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hc)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h2d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h5)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h33: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h46)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h39: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h23)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h3f: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub00_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub01_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub02_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub03_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub04_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub05_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub06_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub07_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sys_run_step <= 7'h0;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= ((w_sub08_run_busy) ? r_sys_run_step : w_sys_run_step_p1);

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h42: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h3a)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h48: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h1d)) begin
										r_sys_run_step <= w_sys_run_step_p1;

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sys_run_step <= 7'h0;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sys_run_busy <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h0: begin
					r_sys_run_busy <= ((i_run_req) ? w_sys_boolTrue : w_sys_boolFalse);
				end

				2'h1: begin

					case(r_sys_run_phase) 
						7'h0: begin
							r_sys_run_busy <= w_sys_boolTrue;
						end

						7'h4d: begin
							r_sys_run_busy <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp23[8:0] );

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1485[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1489[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1481[8:0] );

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1503[8:0] );

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h2) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1498[8:0] );

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1589[8:0] );

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1845[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1953[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1803[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1647[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1809[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1833[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2007[8:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2031[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1641[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1731[8:0] );

									end
									else
									if((r_sys_run_step==7'h39) || (r_sys_run_step==7'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1977[8:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2037[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1665[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1755[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1635[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1683[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1851[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1761[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1677[8:0] );

									end
									else
									if((r_sys_run_step==7'h17) || (r_sys_run_step==7'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1773[8:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2019[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1653[8:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2049[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1983[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2013[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1821[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1881[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1971[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1695[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1887[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1725[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1947[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1659[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1965[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1905[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1959[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1797[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2043[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1749[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1767[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1875[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1839[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1893[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1689[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1791[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1743[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1671[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1815[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1941[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1701[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1857[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1869[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1929[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1737[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1935[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1827[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2001[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e) || (r_sys_run_step==7'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1911[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2025[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1899[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1719[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp1863[8:0] );

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2115[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2067[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2103[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2061[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2229[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2091[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2169[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2241[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2157[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2121[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2181[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2085[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2175[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2127[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2073[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2109[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2145[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2235[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2079[8:0] );

									end
									else
									if((r_sys_run_step==7'h17) || (r_sys_run_step==7'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2199[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2193[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2259[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2223[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2253[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2187[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2163[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2151[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2097[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2217[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2247[8:0] );

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h26)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2461[8:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2506[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2283[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2381[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2401[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2376[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2277[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2486[8:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2511[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2476[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2366[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2271[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2371[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2466[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2531[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2411[8:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2386[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2501[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2313[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2396[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2361[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2319[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2346[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2406[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2441[8:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2556[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2521[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2295[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2456[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2426[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2481[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2516[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2491[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2325[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2541[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2546[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2536[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2436[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2446[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2561[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2496[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2336[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2391[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2471[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2416[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2351[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2289[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2307[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2331[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2526[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2421[8:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2566[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2301[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2451[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2431[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2356[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2341[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2551[8:0] );

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2727[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2589[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2613[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2577[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2601[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2607[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2662[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2717[8:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2631[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2583[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2652[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2647[8:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2687[8:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2692[8:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2625[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2619[8:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2642[8:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2637[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2657[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2722[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2677[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2682[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2672[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2707[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2595[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2697[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2702[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2667[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_T_0_addr_1 <= $signed( w_sys_tmp2712[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp1488;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp1483;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp1501;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp1592;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp38_float;

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp29_float;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp37_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp3_float;

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp34_float;

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp35_float;

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp42_float;

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp41_float;

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp1_float;

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp46_float;

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp27_float;

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp30_float;

									end
									else
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2273;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp0_float;

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp25_float;

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp28_float;

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp39_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp36_float;

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp44_float;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp40_float;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp33_float;

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp45_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp32_float;

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp47_float;

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp2_float;

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp43_float;

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp31_float;

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp26_float;

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp24_float;

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp14_float;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1c)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp11_float;

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp15_float;

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp9_float;

									end
									else
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hb)) begin
										r_fld_T_0_datain_1 <= w_sys_tmp2579;

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp10_float;

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp23_float;

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp18_float;

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp20_float;

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp8_float;

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp5_float;

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp17_float;

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp13_float;

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp16_float;

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp21_float;

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp19_float;

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp12_float;

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp6_float;

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp22_float;

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp7_float;

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_T_0_datain_1 <= r_sys_tmp14_float;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_T_0_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h3)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h45)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h21)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h3b)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'h1e)) begin
										r_fld_T_0_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_T_0_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_TT_1_addr_1 <= $signed( w_sys_tmp28[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_TT_1_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_TT_1_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_TT_1_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_TT_1_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp33[8:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h45)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1060[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp688[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp868[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp664[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp976[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp736[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp568[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp592[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp484[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp628[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp328[8:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1000[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp844[8:0] );

									end
									else
									if((r_sys_run_step==7'h17) || (r_sys_run_step==7'h19)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp508[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp316[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp256[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp556[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp616[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp772[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp820[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp340[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp724[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp928[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp472[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp604[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp424[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp832[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp436[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e) || (r_sys_run_step==7'h30)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp784[8:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1036[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp244[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp676[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp640[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp712[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp412[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp700[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp904[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp988[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp268[8:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1024[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp460[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp544[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp652[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp304[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp856[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h18)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp496[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp280[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp232[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp892[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp400[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp964[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1012[8:0] );

									end
									else
									if((r_sys_run_step==7'h39) || (r_sys_run_step==7'h3b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp916[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp352[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1048[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp880[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp748[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp448[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp760[8:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h10)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1270[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1366[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1402[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1294[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1102[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1126[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1414[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1330[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1162[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1150[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1390[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1282[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1318[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1198[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1114[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1210[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1450[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1174[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1090[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1246[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1258[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1186[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1426[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1462[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1438[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1342[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1138[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1078[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1378[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_U_2_addr_1 <= $signed( w_sys_tmp1306[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_U_2_datain_1 <= w_sys_tmp19;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_U_2_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h45)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_U_2_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_U_2_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_addr_1 <= 9'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp42[8:0] );

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h45)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1060[8:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp688[8:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp868[8:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp664[8:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp976[8:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp736[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp568[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp592[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp484[8:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp628[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp328[8:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1000[8:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp844[8:0] );

									end
									else
									if((r_sys_run_step==7'h17) || (r_sys_run_step==7'h19)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp508[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp316[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp256[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp556[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp616[8:0] );

									end
									else
									if((r_sys_run_step==7'h2d) || (r_sys_run_step==7'h2f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp772[8:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp820[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp340[8:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp724[8:0] );

									end
									else
									if((r_sys_run_step==7'h3a) || (r_sys_run_step==7'h3c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp928[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp472[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp604[8:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp424[8:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp832[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp436[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp364[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp580[8:0] );

									end
									else
									if((r_sys_run_step==7'h2e) || (r_sys_run_step==7'h30)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp784[8:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1036[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp244[8:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp676[8:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp640[8:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp712[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp412[8:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp700[8:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp904[8:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp988[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp268[8:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1024[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp460[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp544[8:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp652[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp304[8:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp856[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h18)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp496[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp280[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp232[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp292[8:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp892[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp400[8:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp964[8:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1012[8:0] );

									end
									else
									if((r_sys_run_step==7'h39) || (r_sys_run_step==7'h3b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp916[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp352[8:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1048[8:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp880[8:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp748[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp448[8:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp760[8:0] );

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h10)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1270[8:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1366[8:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1402[8:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1294[8:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1102[8:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1126[8:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1414[8:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1330[8:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1162[8:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1150[8:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1390[8:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1282[8:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1318[8:0] );

									end
									else
									if((r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1198[8:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1114[8:0] );

									end
									else
									if((r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1210[8:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1450[8:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1174[8:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1090[8:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1246[8:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1258[8:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1186[8:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1426[8:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1462[8:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1438[8:0] );

									end
									else
									if((r_sys_run_step==7'h16) || (r_sys_run_step==7'h17)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1342[8:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1138[8:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1078[8:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1378[8:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_fld_V_3_addr_1 <= $signed( w_sys_tmp1306[8:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_datain_1 <= w_sys_tmp26;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_fld_V_3_r_w_1 <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h45)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_fld_V_3_r_w_1 <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_fld_V_3_r_w_1 <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_13 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h6: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_13 <= w_sys_tmp15;

									end
								end

							endcase
						end

						7'hf: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_13 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_run_k_13 <= w_sys_tmp1071;

									end
								end

							endcase
						end

						7'h15: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_13 <= w_sys_tmp1072;

									end
								end

							endcase
						end

						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h22)) begin
										r_run_k_13 <= w_sys_tmp1473;

									end
								end

							endcase
						end

						7'h20: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_13 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h24: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_run_k_13 <= w_sys_tmp1493;

									end
								end

							endcase
						end

						7'h32: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_13 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_run_k_13 <= w_sys_tmp2054;

									end
								end

							endcase
						end

						7'h38: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_13 <= w_sys_tmp2055;

									end
								end

							endcase
						end

						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h23)) begin
										r_run_k_13 <= w_sys_tmp2264;

									end
								end

							endcase
						end

						7'h41: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_13 <= w_sys_tmp2265;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3b)) begin
										r_run_k_13 <= w_sys_tmp2570;

									end
								end

							endcase
						end

						7'h47: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_k_13 <= w_sys_tmp2571;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_run_k_13 <= w_sys_tmp2731;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_14 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_14 <= w_sys_tmp49;

									end
								end

							endcase
						end

						7'h26: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_14 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0) || (r_sys_run_step==7'h2) || (r_sys_run_step==7'h4) || (r_sys_run_step==7'h6) || (r_sys_run_step==7'h8) || (r_sys_run_step==7'ha) || (r_sys_run_step==7'hc)) begin
										r_run_j_14 <= w_sys_tmp1508;

									end
								end

							endcase
						end

						7'h2c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_j_14 <= w_sys_tmp1581;

									end
								end

							endcase
						end

						7'h30: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_j_14 <= w_sys_tmp1593;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h1b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_15 <= w_sys_intOne;

									end
								end

							endcase
						end

						7'h1d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_n_15 <= w_sys_tmp1476;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_mx_16 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_my_17 <= w_sys_tmp3;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dt_18 <= w_sys_tmp5;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dx_19 <= w_sys_tmp7;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_dy_20 <= w_sys_tmp8;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r1_21 <= w_sys_tmp9;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r2_22 <= w_sys_tmp10;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r3_23 <= w_sys_tmp11;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_r4_24 <= w_sys_tmp12;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h10) || (r_sys_run_step==7'h11)) begin
										r_run_YY_25 <= r_sys_tmp4_float;

									end
									else
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'hd) || (r_sys_run_step==7'he) || (r_sys_run_step==7'h12) || (r_sys_run_step==7'h14)) begin
										r_run_YY_25 <= w_sys_tmp19;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_kx_26 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_ky_27 <= w_sys_tmp1;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h2: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_nlast_28 <= w_sys_tmp6;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_29 <= r_run_j_14;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy0_j_29 <= w_sys_tmp46;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy1_j_30 <= r_run_j_14;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h18) || (r_sys_run_step==7'h1a) || (7'h1c<=r_sys_run_step && r_sys_run_step<=7'h20)) begin
										r_run_copy1_j_30 <= w_sys_tmp47;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h9: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy2_j_31 <= r_run_j_14;

									end
								end

							endcase
						end

						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h6)) begin
										r_run_copy2_j_31 <= w_sys_tmp48;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h26: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_run_copy0_j_32 <= r_run_j_14;

									end
								end

							endcase
						end

						7'h2a: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1) || (r_sys_run_step==7'h3) || (r_sys_run_step==7'h5) || (r_sys_run_step==7'h7) || (r_sys_run_step==7'h9) || (r_sys_run_step==7'hb) || (r_sys_run_step==7'hd)) begin
										r_run_copy0_j_32 <= w_sys_tmp1507;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h8: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub08_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub08_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1d)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2223[9:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2253[9:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2241[9:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2235[9:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2199[9:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2193[9:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2229[9:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2217[9:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2247[9:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_sub08_T_addr <= $signed( w_sys_tmp2259[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h23)) begin
										r_sub08_T_datain <= w_sys_tmp2063;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h23)) begin
										r_sub08_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h21)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1450[9:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1414[9:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1366[9:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1462[9:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1402[9:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1438[9:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1342[9:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1390[9:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1378[9:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub08_V_addr <= $signed( w_sys_tmp1426[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub08_V_datain <= w_sys_tmp1086;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub08_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h21)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1450[9:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1414[9:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1366[9:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1462[9:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1402[9:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1438[9:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1342[9:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1390[9:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1378[9:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub08_U_addr <= $signed( w_sys_tmp1426[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub08_U_datain <= w_sys_tmp1080;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h19<=r_sys_run_step && r_sys_run_step<=7'h22)) begin
										r_sub08_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2707[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2697[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2727[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2717[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2702[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2722[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2712[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2687[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub08_result_addr <= $signed( w_sys_tmp2692[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub08_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub08_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub08_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h3: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub03_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h25)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1845[9:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1893[9:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1869[9:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1905[9:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1875[9:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1851[9:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1881[9:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1911[9:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1887[9:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1899[9:0] );

									end
									else
									if((r_sys_run_step==7'h28)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1863[9:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_sub03_T_addr <= $signed( w_sys_tmp1857[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h25<=r_sys_run_step && r_sys_run_step<=7'h30)) begin
										r_sub03_T_datain <= w_sys_tmp1637;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h25<=r_sys_run_step && r_sys_run_step<=7'h30)) begin
										r_sub03_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h28)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp688[9:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp784[9:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp724[9:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp748[9:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp676[9:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp664[9:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp772[9:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp652[9:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp736[9:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp712[9:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp760[9:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_sub03_V_addr <= $signed( w_sys_tmp700[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h25<=r_sys_run_step && r_sys_run_step<=7'h30)) begin
										r_sub03_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h25<=r_sys_run_step && r_sys_run_step<=7'h30)) begin
										r_sub03_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h28)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp688[9:0] );

									end
									else
									if((r_sys_run_step==7'h30)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp784[9:0] );

									end
									else
									if((r_sys_run_step==7'h2b)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp724[9:0] );

									end
									else
									if((r_sys_run_step==7'h2d)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp748[9:0] );

									end
									else
									if((r_sys_run_step==7'h27)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp676[9:0] );

									end
									else
									if((r_sys_run_step==7'h26)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp664[9:0] );

									end
									else
									if((r_sys_run_step==7'h2f)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp772[9:0] );

									end
									else
									if((r_sys_run_step==7'h25)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp652[9:0] );

									end
									else
									if((r_sys_run_step==7'h2c)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp736[9:0] );

									end
									else
									if((r_sys_run_step==7'h2a)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp712[9:0] );

									end
									else
									if((r_sys_run_step==7'h2e)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp760[9:0] );

									end
									else
									if((r_sys_run_step==7'h29)) begin
										r_sub03_U_addr <= $signed( w_sys_tmp700[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h25<=r_sys_run_step && r_sys_run_step<=7'h30)) begin
										r_sub03_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h25<=r_sys_run_step && r_sys_run_step<=7'h30)) begin
										r_sub03_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2461[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2471[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2466[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2436[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2431[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2456[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2446[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2441[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2426[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub03_result_addr <= $signed( w_sys_tmp2451[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub03_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub03_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub03_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h2: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub02_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub02_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1b)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1773[9:0] );

									end
									else
									if((r_sys_run_step==7'h1e)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1803[9:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1797[9:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1791[9:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1833[9:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1809[9:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1767[9:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1815[9:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1827[9:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1839[9:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub02_T_addr <= $signed( w_sys_tmp1821[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sub02_T_datain <= w_sys_tmp1637;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sub02_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp568[9:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp496[9:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp556[9:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp592[9:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp580[9:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp616[9:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp628[9:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp544[9:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp640[9:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp508[9:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub02_V_addr <= $signed( w_sys_tmp604[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sub02_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sub02_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1e)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp568[9:0] );

									end
									else
									if((r_sys_run_step==7'h1a)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp496[9:0] );

									end
									else
									if((r_sys_run_step==7'h1d)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp556[9:0] );

									end
									else
									if((r_sys_run_step==7'h20)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp592[9:0] );

									end
									else
									if((r_sys_run_step==7'h1f)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp580[9:0] );

									end
									else
									if((r_sys_run_step==7'h22)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp616[9:0] );

									end
									else
									if((r_sys_run_step==7'h23)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp628[9:0] );

									end
									else
									if((r_sys_run_step==7'h1c)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp544[9:0] );

									end
									else
									if((r_sys_run_step==7'h24)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp640[9:0] );

									end
									else
									if((r_sys_run_step==7'h1b)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp508[9:0] );

									end
									else
									if((r_sys_run_step==7'h21)) begin
										r_sub02_U_addr <= $signed( w_sys_tmp604[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sub02_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h1a<=r_sys_run_step && r_sys_run_step<=7'h24)) begin
										r_sub02_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2401[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2381[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2391[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2396[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2411[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2421[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2416[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2406[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub02_result_addr <= $signed( w_sys_tmp2386[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub02_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub02_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub02_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h1: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub01_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub01_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h19)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1773[9:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1737[9:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1767[9:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1743[9:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1761[9:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1755[9:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1695[9:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1731[9:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1725[9:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1749[9:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1719[9:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub01_T_addr <= $signed( w_sys_tmp1701[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub01_T_datain <= w_sys_tmp1637;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub01_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h18)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp496[9:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp436[9:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp364[9:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp472[9:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp400[9:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp484[9:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp460[9:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp448[9:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp508[9:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp352[9:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp412[9:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub01_V_addr <= $signed( w_sys_tmp424[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub01_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub01_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h18)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp496[9:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp436[9:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp364[9:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp472[9:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp400[9:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp484[9:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp460[9:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp448[9:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp508[9:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp352[9:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp412[9:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub01_U_addr <= $signed( w_sys_tmp424[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub01_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub01_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2331[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2366[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2336[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2376[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2371[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2361[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2351[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2356[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2346[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub01_result_addr <= $signed( w_sys_tmp2341[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub01_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub01_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub01_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub00_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub00_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1659[9:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1689[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1653[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1635[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1683[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1671[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1665[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1647[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1677[9:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1695[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1641[9:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub00_T_addr <= $signed( w_sys_tmp1701[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub00_T_datain <= w_sys_tmp1637;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub00_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp364[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp280[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp256[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp232[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp268[9:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp340[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp292[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp244[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp328[9:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp352[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp316[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub00_V_addr <= $signed( w_sys_tmp304[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub00_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub00_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hd)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp364[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp280[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp256[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp232[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp268[9:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp340[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp292[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp244[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp328[9:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp352[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp316[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub00_U_addr <= $signed( w_sys_tmp304[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub00_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub00_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2325[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2307[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2295[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2283[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2313[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2271[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2319[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2277[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2301[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub00_result_addr <= $signed( w_sys_tmp2289[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub00_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub00_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub00_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h7: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub07_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub07_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h14)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2169[9:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2187[9:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2163[9:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2145[9:0] );

									end
									else
									if((r_sys_run_step==7'h19)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2199[9:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2193[9:0] );

									end
									else
									if((r_sys_run_step==7'h12)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2157[9:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2151[9:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2181[9:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2121[9:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2175[9:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub07_T_addr <= $signed( w_sys_tmp2127[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub07_T_datain <= w_sys_tmp2063;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h19)) begin
										r_sub07_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h12)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1270[9:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1198[9:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1210[9:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1330[9:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1342[9:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1246[9:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1294[9:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1282[9:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1258[9:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1318[9:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub07_V_addr <= $signed( w_sys_tmp1306[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub07_V_datain <= w_sys_tmp1086;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub07_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h12)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1270[9:0] );

									end
									else
									if((r_sys_run_step==7'he)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1198[9:0] );

									end
									else
									if((r_sys_run_step==7'hf)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1210[9:0] );

									end
									else
									if((r_sys_run_step==7'h17)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1330[9:0] );

									end
									else
									if((r_sys_run_step==7'h18)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1342[9:0] );

									end
									else
									if((r_sys_run_step==7'h10)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1246[9:0] );

									end
									else
									if((r_sys_run_step==7'h14)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1294[9:0] );

									end
									else
									if((r_sys_run_step==7'h13)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1282[9:0] );

									end
									else
									if((r_sys_run_step==7'h11)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1258[9:0] );

									end
									else
									if((r_sys_run_step==7'h16)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1318[9:0] );

									end
									else
									if((r_sys_run_step==7'h15)) begin
										r_sub07_U_addr <= $signed( w_sys_tmp1306[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub07_U_datain <= w_sys_tmp1080;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'he<=r_sys_run_step && r_sys_run_step<=7'h18)) begin
										r_sub07_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2662[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2642[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2637[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2657[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2682[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2677[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2667[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2652[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2647[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub07_result_addr <= $signed( w_sys_tmp2672[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub07_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub07_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub07_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h6: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub06_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub06_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2115[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2073[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2067[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2109[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2103[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2079[9:0] );

									end
									else
									if((r_sys_run_step==7'hc)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2121[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2061[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2097[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2085[9:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2127[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub06_T_addr <= $signed( w_sys_tmp2091[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub06_T_datain <= w_sys_tmp2063;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3c: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub06_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hc)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1198[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1114[9:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1210[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1126[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1162[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1174[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1090[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1150[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1138[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1078[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1102[9:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub06_V_addr <= $signed( w_sys_tmp1186[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub06_V_datain <= w_sys_tmp1086;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub06_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hc)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1198[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1114[9:0] );

									end
									else
									if((r_sys_run_step==7'hd)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1210[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1126[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1162[9:0] );

									end
									else
									if((r_sys_run_step==7'ha)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1174[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1090[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1150[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1138[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1078[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1102[9:0] );

									end
									else
									if((r_sys_run_step==7'hb)) begin
										r_sub06_U_addr <= $signed( w_sys_tmp1186[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub06_U_datain <= w_sys_tmp1080;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h19: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h2<=r_sys_run_step && r_sys_run_step<=7'hd)) begin
										r_sub06_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2607[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2595[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2631[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2583[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2589[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2613[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2577[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2625[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2619[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub06_result_addr <= $signed( w_sys_tmp2601[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub06_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub06_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub06_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h5: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub05_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub05_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h42)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2019[9:0] );

									end
									else
									if((r_sys_run_step==7'h47)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2049[9:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp1983[9:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2037[9:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2013[9:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2007[9:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2031[9:0] );

									end
									else
									if((r_sys_run_step==7'h46)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2043[9:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2001[9:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp2025[9:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_sub05_T_addr <= $signed( w_sys_tmp1977[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h3d<=r_sys_run_step && r_sys_run_step<=7'h47)) begin
										r_sub05_T_datain <= w_sys_tmp1637;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h3d<=r_sys_run_step && r_sys_run_step<=7'h47)) begin
										r_sub05_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1060[9:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp988[9:0] );

									end
									else
									if((r_sys_run_step==7'h46)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1048[9:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp928[9:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1036[9:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp964[9:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1024[9:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp976[9:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1012[9:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp916[9:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_sub05_V_addr <= $signed( w_sys_tmp1000[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h3d<=r_sys_run_step && r_sys_run_step<=7'h47)) begin
										r_sub05_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h3d<=r_sys_run_step && r_sys_run_step<=7'h47)) begin
										r_sub05_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h47)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1060[9:0] );

									end
									else
									if((r_sys_run_step==7'h41)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp988[9:0] );

									end
									else
									if((r_sys_run_step==7'h46)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1048[9:0] );

									end
									else
									if((r_sys_run_step==7'h3e)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp928[9:0] );

									end
									else
									if((r_sys_run_step==7'h45)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1036[9:0] );

									end
									else
									if((r_sys_run_step==7'h3f)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp964[9:0] );

									end
									else
									if((r_sys_run_step==7'h44)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1024[9:0] );

									end
									else
									if((r_sys_run_step==7'h40)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp976[9:0] );

									end
									else
									if((r_sys_run_step==7'h43)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1012[9:0] );

									end
									else
									if((r_sys_run_step==7'h3d)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp916[9:0] );

									end
									else
									if((r_sys_run_step==7'h42)) begin
										r_sub05_U_addr <= $signed( w_sys_tmp1000[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h3d<=r_sys_run_step && r_sys_run_step<=7'h47)) begin
										r_sub05_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h3d<=r_sys_run_step && r_sys_run_step<=7'h47)) begin
										r_sub05_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2541[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2526[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2546[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2536[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2531[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2566[9:0] );

									end
									else
									if((r_sys_run_step==7'h6)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2556[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2551[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub05_result_addr <= $signed( w_sys_tmp2561[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub05_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h8)) begin
										r_sub05_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub05_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_run_req <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h4: begin
									if((r_sys_run_step==7'h1)) begin
										r_sub04_run_req <= w_sys_boolFalse;

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub04_run_req <= w_sys_boolTrue;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h36)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1947[9:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1953[9:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1929[9:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1965[9:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1905[9:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1959[9:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1983[9:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1935[9:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1941[9:0] );

									end
									else
									if((r_sys_run_step==7'h3a)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1971[9:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1911[9:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sub04_T_addr <= $signed( w_sys_tmp1977[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h31<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sub04_T_datain <= w_sys_tmp1637;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_T_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h36: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h31<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sub04_T_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_T_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_T_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3a)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp904[9:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp868[9:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp784[9:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp928[9:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp892[9:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp880[9:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp772[9:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp916[9:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp844[9:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp820[9:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp856[9:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_sub04_V_addr <= $signed( w_sys_tmp832[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h31<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sub04_V_datain <= w_sys_tmp240;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_V_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h31<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sub04_V_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_V_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_V_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3a)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp904[9:0] );

									end
									else
									if((r_sys_run_step==7'h37)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp868[9:0] );

									end
									else
									if((r_sys_run_step==7'h32)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp784[9:0] );

									end
									else
									if((r_sys_run_step==7'h3c)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp928[9:0] );

									end
									else
									if((r_sys_run_step==7'h39)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp892[9:0] );

									end
									else
									if((r_sys_run_step==7'h38)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp880[9:0] );

									end
									else
									if((r_sys_run_step==7'h31)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp772[9:0] );

									end
									else
									if((r_sys_run_step==7'h3b)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp916[9:0] );

									end
									else
									if((r_sys_run_step==7'h35)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp844[9:0] );

									end
									else
									if((r_sys_run_step==7'h33)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp820[9:0] );

									end
									else
									if((r_sys_run_step==7'h36)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp856[9:0] );

									end
									else
									if((r_sys_run_step==7'h34)) begin
										r_sub04_U_addr <= $signed( w_sys_tmp832[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h31<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sub04_U_datain <= w_sys_tmp234;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_U_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h13: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h31<=r_sys_run_step && r_sys_run_step<=7'h3c)) begin
										r_sub04_U_r_w <= w_sys_boolTrue;

									end
								end

							endcase
						end

						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_U_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_U_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_addr <= 10'sh0;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2506[9:0] );

									end
									else
									if((r_sys_run_step==7'h5)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2501[9:0] );

									end
									else
									if((r_sys_run_step==7'h4)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2496[9:0] );

									end
									else
									if((r_sys_run_step==7'h7)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2511[9:0] );

									end
									else
									if((r_sys_run_step==7'h2)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2486[9:0] );

									end
									else
									if((r_sys_run_step==7'h8)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2516[9:0] );

									end
									else
									if((r_sys_run_step==7'h1)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2481[9:0] );

									end
									else
									if((r_sys_run_step==7'h9)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2521[9:0] );

									end
									else
									if((r_sys_run_step==7'h3)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2491[9:0] );

									end
									else
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_addr <= $signed( w_sys_tmp2476[9:0] );

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(( !reset_n )) begin
			r_sub04_result_r_w <= w_sys_boolFalse;

		end
		else
		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h3d: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h1: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h2: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h3: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h4: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h5: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h6: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h7: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

								4'h8: begin
									if((r_sys_run_step==7'h0)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((7'h0<=r_sys_run_step && r_sys_run_step<=7'h9)) begin
										r_sub04_result_r_w <= w_sys_boolFalse;

									end
								end

							endcase
						end

						7'h4d: begin
							r_sub04_result_r_w <= w_sys_boolFalse;
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_tmp0_float <= w_ip_MultFloat_product_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp0_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h16)) begin
										r_sys_tmp1_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp1_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h12) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h19)) begin
										r_sys_tmp2_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp2_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h17)) begin
										r_sys_tmp3_float <= w_ip_AddFloat_result_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp3_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'hd: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hf) || (r_sys_run_step==7'h10) || (r_sys_run_step==7'h11) || (r_sys_run_step==7'h13) || (r_sys_run_step==7'h15) || (r_sys_run_step==7'h17) || (r_sys_run_step==7'h19)) begin
										r_sys_tmp4_float <= w_ip_MultFloat_product_0;

									end
									else
									if((r_sys_run_step==7'hc) || (r_sys_run_step==7'hd)) begin
										r_sys_tmp4_float <= w_ip_FixedToFloat_floating_0;

									end
								end

							endcase
						end

						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp4_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp5_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'hb)) begin
										r_sys_tmp5_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp6_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp6_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp7_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'ha)) begin
										r_sys_tmp7_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp8_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp8_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp9_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp9_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp10_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp10_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp11_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp11_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h9)) begin
										r_sys_tmp12_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp12_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp13_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp13_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp14_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp14_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp15_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp15_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp16_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp16_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h8)) begin
										r_sys_tmp17_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp17_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp18_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp18_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp19_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp19_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp20_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp20_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp21_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp21_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h7)) begin
										r_sys_tmp22_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp22_float <= w_sub08_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp23_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

						7'h4b: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp23_float <= w_sub07_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp24_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp25_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp26_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h6)) begin
										r_sys_tmp27_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp28_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp29_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp30_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp31_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h5)) begin
										r_sys_tmp32_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp33_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp34_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp35_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp36_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h4)) begin
										r_sys_tmp37_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp38_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp39_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp40_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp41_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h3)) begin
										r_sys_tmp42_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp43_float <= w_sub01_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp44_float <= w_sub04_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp45_float <= w_sub03_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp46_float <= w_sub05_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


	always@(posedge clock)begin

		if(w_sys_ce) begin

			case(r_sys_processing_methodID) 
				2'h1: begin

					case(r_sys_run_phase) 
						7'h45: begin

							case(r_sys_run_stage) 
								4'h0: begin
									if((r_sys_run_step==7'h2)) begin
										r_sys_tmp47_float <= w_sub02_result_dataout;

									end
								end

							endcase
						end

					endcase
				end

			endcase
		end
	end


endmodule
